

module padder53(A, B, Cin, S, Cout);
  parameter N = 53;
  input [N-1:0] A, B;
  input Cin;
  output [N-1:0] S;
  output Cout;

  // P[i] is an alias for Pi:i, likewise G[i] is an alias for Gi:i
  wire [N-2:-1] P, G;

  assign P = {A[N-2:0] | B[N-2:0], 1'b0};
  assign G = {A[N-2:0] & B[N-2:0], Cin};

  Sum s0(G[-1], A[0], B[0], S[0]);

  wire \G0:-1 ;

  Gij \0:-1 (P[0], G[0], G[-1], \G0:-1 );

  Sum s1(\G0:-1 , A[1], B[1], S[1]);

  wire \G1:-1 ;

  Gij \1:-1 (P[1], G[1], \G0:-1 , \G1:-1 );

  Sum s2(\G1:-1 , A[2], B[2], S[2]);

  wire \P2:1 , \G2:1 ;

  PijGij \2:1 (P[2], P[1], G[2], G[1], \P2:1 , \G2:1 );

  wire \G2:-1 ;

  Gij \2:-1 (\P2:1 , \G2:1 , \G0:-1 , \G2:-1 );

  Sum s3(\G2:-1 , A[3], B[3], S[3]);

  wire \G3:-1 ;

  Gij \3:-1 (P[3], G[3], \G2:-1 , \G3:-1 );

  Sum s4(\G3:-1 , A[4], B[4], S[4]);

  wire \P4:3 , \G4:3 ;

  PijGij \4:3 (P[4], P[3], G[4], G[3], \P4:3 , \G4:3 );

  wire \G4:-1 ;

  Gij \4:-1 (\P4:3 , \G4:3 , \G2:-1 , \G4:-1 );

  Sum s5(\G4:-1 , A[5], B[5], S[5]);

  wire \P5:3 , \G5:3 ;

  PijGij \5:3 (P[5], \P4:3 , G[5], \G4:3 , \P5:3 , \G5:3 );

  wire \G5:-1 ;

  Gij \5:-1 (\P5:3 , \G5:3 , \G2:-1 , \G5:-1 );

  Sum s6(\G5:-1 , A[6], B[6], S[6]);

  wire \P6:5 , \G6:5 ;

  PijGij \6:5 (P[6], P[5], G[6], G[5], \P6:5 , \G6:5 );

  wire \P6:3 , \G6:3 ;

  PijGij \6:3 (\P6:5 , \P4:3 , \G6:5 , \G4:3 , \P6:3 , \G6:3 );

  wire \G6:-1 ;

  Gij \6:-1 (\P6:3 , \G6:3 , \G2:-1 , \G6:-1 );

  Sum s7(\G6:-1 , A[7], B[7], S[7]);

  wire \G7:-1 ;

  Gij \7:-1 (P[7], G[7], \G6:-1 , \G7:-1 );

  Sum s8(\G7:-1 , A[8], B[8], S[8]);

  wire \P8:7 , \G8:7 ;

  PijGij \8:7 (P[8], P[7], G[8], G[7], \P8:7 , \G8:7 );

  wire \G8:-1 ;

  Gij \8:-1 (\P8:7 , \G8:7 , \G6:-1 , \G8:-1 );

  Sum s9(\G8:-1 , A[9], B[9], S[9]);

  wire \P9:7 , \G9:7 ;

  PijGij \9:7 (P[9], \P8:7 , G[9], \G8:7 , \P9:7 , \G9:7 );

  wire \G9:-1 ;

  Gij \9:-1 (\P9:7 , \G9:7 , \G6:-1 , \G9:-1 );

  Sum s10(\G9:-1 , A[10], B[10], S[10]);

  wire \P10:9 , \G10:9 ;

  PijGij \10:9 (P[10], P[9], G[10], G[9], \P10:9 , \G10:9 );

  wire \P10:7 , \G10:7 ;

  PijGij \10:7 (\P10:9 , \P8:7 , \G10:9 , \G8:7 , \P10:7 , \G10:7 );

  wire \G10:-1 ;

  Gij \10:-1 (\P10:7 , \G10:7 , \G6:-1 , \G10:-1 );

  Sum s11(\G10:-1 , A[11], B[11], S[11]);

  wire \P11:7 , \G11:7 ;

  PijGij \11:7 (P[11], \P10:7 , G[11], \G10:7 , \P11:7 , \G11:7 );

  wire \G11:-1 ;

  Gij \11:-1 (\P11:7 , \G11:7 , \G6:-1 , \G11:-1 );

  Sum s12(\G11:-1 , A[12], B[12], S[12]);

  wire \P12:11 , \G12:11 ;

  PijGij \12:11 (P[12], P[11], G[12], G[11], \P12:11 , \G12:11 );

  wire \P12:7 , \G12:7 ;

  PijGij \12:7 (\P12:11 , \P10:7 , \G12:11 , \G10:7 , \P12:7 , \G12:7 );

  wire \G12:-1 ;

  Gij \12:-1 (\P12:7 , \G12:7 , \G6:-1 , \G12:-1 );

  Sum s13(\G12:-1 , A[13], B[13], S[13]);

  wire \P13:11 , \G13:11 ;

  PijGij \13:11 (P[13], \P12:11 , G[13], \G12:11 , \P13:11 , \G13:11 );

  wire \P13:7 , \G13:7 ;

  PijGij \13:7 (\P13:11 , \P10:7 , \G13:11 , \G10:7 , \P13:7 , \G13:7 );

  wire \G13:-1 ;

  Gij \13:-1 (\P13:7 , \G13:7 , \G6:-1 , \G13:-1 );

  Sum s14(\G13:-1 , A[14], B[14], S[14]);

  wire \P14:13 , \G14:13 ;

  PijGij \14:13 (P[14], P[13], G[14], G[13], \P14:13 , \G14:13 );

  wire \P14:11 , \G14:11 ;

  PijGij \14:11 (\P14:13 , \P12:11 , \G14:13 , \G12:11 , \P14:11 , \G14:11 );

  wire \P14:7 , \G14:7 ;

  PijGij \14:7 (\P14:11 , \P10:7 , \G14:11 , \G10:7 , \P14:7 , \G14:7 );

  wire \G14:-1 ;

  Gij \14:-1 (\P14:7 , \G14:7 , \G6:-1 , \G14:-1 );

  Sum s15(\G14:-1 , A[15], B[15], S[15]);

  wire \G15:-1 ;

  Gij \15:-1 (P[15], G[15], \G14:-1 , \G15:-1 );

  Sum s16(\G15:-1 , A[16], B[16], S[16]);

  wire \P16:15 , \G16:15 ;

  PijGij \16:15 (P[16], P[15], G[16], G[15], \P16:15 , \G16:15 );

  wire \G16:-1 ;

  Gij \16:-1 (\P16:15 , \G16:15 , \G14:-1 , \G16:-1 );

  Sum s17(\G16:-1 , A[17], B[17], S[17]);

  wire \P17:15 , \G17:15 ;

  PijGij \17:15 (P[17], \P16:15 , G[17], \G16:15 , \P17:15 , \G17:15 );

  wire \G17:-1 ;

  Gij \17:-1 (\P17:15 , \G17:15 , \G14:-1 , \G17:-1 );

  Sum s18(\G17:-1 , A[18], B[18], S[18]);

  wire \P18:17 , \G18:17 ;

  PijGij \18:17 (P[18], P[17], G[18], G[17], \P18:17 , \G18:17 );

  wire \P18:15 , \G18:15 ;

  PijGij \18:15 (\P18:17 , \P16:15 , \G18:17 , \G16:15 , \P18:15 , \G18:15 );

  wire \G18:-1 ;

  Gij \18:-1 (\P18:15 , \G18:15 , \G14:-1 , \G18:-1 );

  Sum s19(\G18:-1 , A[19], B[19], S[19]);

  wire \P19:15 , \G19:15 ;

  PijGij \19:15 (P[19], \P18:15 , G[19], \G18:15 , \P19:15 , \G19:15 );

  wire \G19:-1 ;

  Gij \19:-1 (\P19:15 , \G19:15 , \G14:-1 , \G19:-1 );

  Sum s20(\G19:-1 , A[20], B[20], S[20]);

  wire \P20:19 , \G20:19 ;

  PijGij \20:19 (P[20], P[19], G[20], G[19], \P20:19 , \G20:19 );

  wire \P20:15 , \G20:15 ;

  PijGij \20:15 (\P20:19 , \P18:15 , \G20:19 , \G18:15 , \P20:15 , \G20:15 );

  wire \G20:-1 ;

  Gij \20:-1 (\P20:15 , \G20:15 , \G14:-1 , \G20:-1 );

  Sum s21(\G20:-1 , A[21], B[21], S[21]);

  wire \P21:19 , \G21:19 ;

  PijGij \21:19 (P[21], \P20:19 , G[21], \G20:19 , \P21:19 , \G21:19 );

  wire \P21:15 , \G21:15 ;

  PijGij \21:15 (\P21:19 , \P18:15 , \G21:19 , \G18:15 , \P21:15 , \G21:15 );

  wire \G21:-1 ;

  Gij \21:-1 (\P21:15 , \G21:15 , \G14:-1 , \G21:-1 );

  Sum s22(\G21:-1 , A[22], B[22], S[22]);

  wire \P22:21 , \G22:21 ;

  PijGij \22:21 (P[22], P[21], G[22], G[21], \P22:21 , \G22:21 );

  wire \P22:19 , \G22:19 ;

  PijGij \22:19 (\P22:21 , \P20:19 , \G22:21 , \G20:19 , \P22:19 , \G22:19 );

  wire \P22:15 , \G22:15 ;

  PijGij \22:15 (\P22:19 , \P18:15 , \G22:19 , \G18:15 , \P22:15 , \G22:15 );

  wire \G22:-1 ;

  Gij \22:-1 (\P22:15 , \G22:15 , \G14:-1 , \G22:-1 );

  Sum s23(\G22:-1 , A[23], B[23], S[23]);

  wire \P23:15 , \G23:15 ;

  PijGij \23:15 (P[23], \P22:15 , G[23], \G22:15 , \P23:15 , \G23:15 );

  wire \G23:-1 ;

  Gij \23:-1 (\P23:15 , \G23:15 , \G14:-1 , \G23:-1 );

  Sum s24(\G23:-1 , A[24], B[24], S[24]);

  wire \P24:23 , \G24:23 ;

  PijGij \24:23 (P[24], P[23], G[24], G[23], \P24:23 , \G24:23 );

  wire \P24:15 , \G24:15 ;

  PijGij \24:15 (\P24:23 , \P22:15 , \G24:23 , \G22:15 , \P24:15 , \G24:15 );

  wire \G24:-1 ;

  Gij \24:-1 (\P24:15 , \G24:15 , \G14:-1 , \G24:-1 );

  Sum s25(\G24:-1 , A[25], B[25], S[25]);

  wire \P25:23 , \G25:23 ;

  PijGij \25:23 (P[25], \P24:23 , G[25], \G24:23 , \P25:23 , \G25:23 );

  wire \P25:15 , \G25:15 ;

  PijGij \25:15 (\P25:23 , \P22:15 , \G25:23 , \G22:15 , \P25:15 , \G25:15 );

  wire \G25:-1 ;

  Gij \25:-1 (\P25:15 , \G25:15 , \G14:-1 , \G25:-1 );

  Sum s26(\G25:-1 , A[26], B[26], S[26]);

  wire \P26:25 , \G26:25 ;

  PijGij \26:25 (P[26], P[25], G[26], G[25], \P26:25 , \G26:25 );

  wire \P26:23 , \G26:23 ;

  PijGij \26:23 (\P26:25 , \P24:23 , \G26:25 , \G24:23 , \P26:23 , \G26:23 );

  wire \P26:15 , \G26:15 ;

  PijGij \26:15 (\P26:23 , \P22:15 , \G26:23 , \G22:15 , \P26:15 , \G26:15 );

  wire \G26:-1 ;

  Gij \26:-1 (\P26:15 , \G26:15 , \G14:-1 , \G26:-1 );

  Sum s27(\G26:-1 , A[27], B[27], S[27]);

  wire \P27:23 , \G27:23 ;

  PijGij \27:23 (P[27], \P26:23 , G[27], \G26:23 , \P27:23 , \G27:23 );

  wire \P27:15 , \G27:15 ;

  PijGij \27:15 (\P27:23 , \P22:15 , \G27:23 , \G22:15 , \P27:15 , \G27:15 );

  wire \G27:-1 ;

  Gij \27:-1 (\P27:15 , \G27:15 , \G14:-1 , \G27:-1 );

  Sum s28(\G27:-1 , A[28], B[28], S[28]);

  wire \P28:27 , \G28:27 ;

  PijGij \28:27 (P[28], P[27], G[28], G[27], \P28:27 , \G28:27 );

  wire \P28:23 , \G28:23 ;

  PijGij \28:23 (\P28:27 , \P26:23 , \G28:27 , \G26:23 , \P28:23 , \G28:23 );

  wire \P28:15 , \G28:15 ;

  PijGij \28:15 (\P28:23 , \P22:15 , \G28:23 , \G22:15 , \P28:15 , \G28:15 );

  wire \G28:-1 ;

  Gij \28:-1 (\P28:15 , \G28:15 , \G14:-1 , \G28:-1 );

  Sum s29(\G28:-1 , A[29], B[29], S[29]);

  wire \P29:27 , \G29:27 ;

  PijGij \29:27 (P[29], \P28:27 , G[29], \G28:27 , \P29:27 , \G29:27 );

  wire \P29:23 , \G29:23 ;

  PijGij \29:23 (\P29:27 , \P26:23 , \G29:27 , \G26:23 , \P29:23 , \G29:23 );

  wire \P29:15 , \G29:15 ;

  PijGij \29:15 (\P29:23 , \P22:15 , \G29:23 , \G22:15 , \P29:15 , \G29:15 );

  wire \G29:-1 ;

  Gij \29:-1 (\P29:15 , \G29:15 , \G14:-1 , \G29:-1 );

  Sum s30(\G29:-1 , A[30], B[30], S[30]);

  wire \P30:29 , \G30:29 ;

  PijGij \30:29 (P[30], P[29], G[30], G[29], \P30:29 , \G30:29 );

  wire \P30:27 , \G30:27 ;

  PijGij \30:27 (\P30:29 , \P28:27 , \G30:29 , \G28:27 , \P30:27 , \G30:27 );

  wire \P30:23 , \G30:23 ;

  PijGij \30:23 (\P30:27 , \P26:23 , \G30:27 , \G26:23 , \P30:23 , \G30:23 );

  wire \P30:15 , \G30:15 ;

  PijGij \30:15 (\P30:23 , \P22:15 , \G30:23 , \G22:15 , \P30:15 , \G30:15 );

  wire \G30:-1 ;

  Gij \30:-1 (\P30:15 , \G30:15 , \G14:-1 , \G30:-1 );

  Sum s31(\G30:-1 , A[31], B[31], S[31]);

  wire \G31:-1 ;

  Gij \31:-1 (P[31], G[31], \G30:-1 , \G31:-1 );

  Sum s32(\G31:-1 , A[32], B[32], S[32]);

  wire \P32:31 , \G32:31 ;

  PijGij \32:31 (P[32], P[31], G[32], G[31], \P32:31 , \G32:31 );

  wire \G32:-1 ;

  Gij \32:-1 (\P32:31 , \G32:31 , \G30:-1 , \G32:-1 );

  Sum s33(\G32:-1 , A[33], B[33], S[33]);

  wire \P33:31 , \G33:31 ;

  PijGij \33:31 (P[33], \P32:31 , G[33], \G32:31 , \P33:31 , \G33:31 );

  wire \G33:-1 ;

  Gij \33:-1 (\P33:31 , \G33:31 , \G30:-1 , \G33:-1 );

  Sum s34(\G33:-1 , A[34], B[34], S[34]);

  wire \P34:33 , \G34:33 ;

  PijGij \34:33 (P[34], P[33], G[34], G[33], \P34:33 , \G34:33 );

  wire \P34:31 , \G34:31 ;

  PijGij \34:31 (\P34:33 , \P32:31 , \G34:33 , \G32:31 , \P34:31 , \G34:31 );

  wire \G34:-1 ;

  Gij \34:-1 (\P34:31 , \G34:31 , \G30:-1 , \G34:-1 );

  Sum s35(\G34:-1 , A[35], B[35], S[35]);

  wire \P35:31 , \G35:31 ;

  PijGij \35:31 (P[35], \P34:31 , G[35], \G34:31 , \P35:31 , \G35:31 );

  wire \G35:-1 ;

  Gij \35:-1 (\P35:31 , \G35:31 , \G30:-1 , \G35:-1 );

  Sum s36(\G35:-1 , A[36], B[36], S[36]);

  wire \P36:35 , \G36:35 ;

  PijGij \36:35 (P[36], P[35], G[36], G[35], \P36:35 , \G36:35 );

  wire \P36:31 , \G36:31 ;

  PijGij \36:31 (\P36:35 , \P34:31 , \G36:35 , \G34:31 , \P36:31 , \G36:31 );

  wire \G36:-1 ;

  Gij \36:-1 (\P36:31 , \G36:31 , \G30:-1 , \G36:-1 );

  Sum s37(\G36:-1 , A[37], B[37], S[37]);

  wire \P37:35 , \G37:35 ;

  PijGij \37:35 (P[37], \P36:35 , G[37], \G36:35 , \P37:35 , \G37:35 );

  wire \P37:31 , \G37:31 ;

  PijGij \37:31 (\P37:35 , \P34:31 , \G37:35 , \G34:31 , \P37:31 , \G37:31 );

  wire \G37:-1 ;

  Gij \37:-1 (\P37:31 , \G37:31 , \G30:-1 , \G37:-1 );

  Sum s38(\G37:-1 , A[38], B[38], S[38]);

  wire \P38:37 , \G38:37 ;

  PijGij \38:37 (P[38], P[37], G[38], G[37], \P38:37 , \G38:37 );

  wire \P38:35 , \G38:35 ;

  PijGij \38:35 (\P38:37 , \P36:35 , \G38:37 , \G36:35 , \P38:35 , \G38:35 );

  wire \P38:31 , \G38:31 ;

  PijGij \38:31 (\P38:35 , \P34:31 , \G38:35 , \G34:31 , \P38:31 , \G38:31 );

  wire \G38:-1 ;

  Gij \38:-1 (\P38:31 , \G38:31 , \G30:-1 , \G38:-1 );

  Sum s39(\G38:-1 , A[39], B[39], S[39]);

  wire \P39:31 , \G39:31 ;

  PijGij \39:31 (P[39], \P38:31 , G[39], \G38:31 , \P39:31 , \G39:31 );

  wire \G39:-1 ;

  Gij \39:-1 (\P39:31 , \G39:31 , \G30:-1 , \G39:-1 );

  Sum s40(\G39:-1 , A[40], B[40], S[40]);

  wire \P40:39 , \G40:39 ;

  PijGij \40:39 (P[40], P[39], G[40], G[39], \P40:39 , \G40:39 );

  wire \P40:31 , \G40:31 ;

  PijGij \40:31 (\P40:39 , \P38:31 , \G40:39 , \G38:31 , \P40:31 , \G40:31 );

  wire \G40:-1 ;

  Gij \40:-1 (\P40:31 , \G40:31 , \G30:-1 , \G40:-1 );

  Sum s41(\G40:-1 , A[41], B[41], S[41]);

  wire \P41:39 , \G41:39 ;

  PijGij \41:39 (P[41], \P40:39 , G[41], \G40:39 , \P41:39 , \G41:39 );

  wire \P41:31 , \G41:31 ;

  PijGij \41:31 (\P41:39 , \P38:31 , \G41:39 , \G38:31 , \P41:31 , \G41:31 );

  wire \G41:-1 ;

  Gij \41:-1 (\P41:31 , \G41:31 , \G30:-1 , \G41:-1 );

  Sum s42(\G41:-1 , A[42], B[42], S[42]);

  wire \P42:41 , \G42:41 ;

  PijGij \42:41 (P[42], P[41], G[42], G[41], \P42:41 , \G42:41 );

  wire \P42:39 , \G42:39 ;

  PijGij \42:39 (\P42:41 , \P40:39 , \G42:41 , \G40:39 , \P42:39 , \G42:39 );

  wire \P42:31 , \G42:31 ;

  PijGij \42:31 (\P42:39 , \P38:31 , \G42:39 , \G38:31 , \P42:31 , \G42:31 );

  wire \G42:-1 ;

  Gij \42:-1 (\P42:31 , \G42:31 , \G30:-1 , \G42:-1 );

  Sum s43(\G42:-1 , A[43], B[43], S[43]);

  wire \P43:39 , \G43:39 ;

  PijGij \43:39 (P[43], \P42:39 , G[43], \G42:39 , \P43:39 , \G43:39 );

  wire \P43:31 , \G43:31 ;

  PijGij \43:31 (\P43:39 , \P38:31 , \G43:39 , \G38:31 , \P43:31 , \G43:31 );

  wire \G43:-1 ;

  Gij \43:-1 (\P43:31 , \G43:31 , \G30:-1 , \G43:-1 );

  Sum s44(\G43:-1 , A[44], B[44], S[44]);

  wire \P44:43 , \G44:43 ;

  PijGij \44:43 (P[44], P[43], G[44], G[43], \P44:43 , \G44:43 );

  wire \P44:39 , \G44:39 ;

  PijGij \44:39 (\P44:43 , \P42:39 , \G44:43 , \G42:39 , \P44:39 , \G44:39 );

  wire \P44:31 , \G44:31 ;

  PijGij \44:31 (\P44:39 , \P38:31 , \G44:39 , \G38:31 , \P44:31 , \G44:31 );

  wire \G44:-1 ;

  Gij \44:-1 (\P44:31 , \G44:31 , \G30:-1 , \G44:-1 );

  Sum s45(\G44:-1 , A[45], B[45], S[45]);

  wire \P45:43 , \G45:43 ;

  PijGij \45:43 (P[45], \P44:43 , G[45], \G44:43 , \P45:43 , \G45:43 );

  wire \P45:39 , \G45:39 ;

  PijGij \45:39 (\P45:43 , \P42:39 , \G45:43 , \G42:39 , \P45:39 , \G45:39 );

  wire \P45:31 , \G45:31 ;

  PijGij \45:31 (\P45:39 , \P38:31 , \G45:39 , \G38:31 , \P45:31 , \G45:31 );

  wire \G45:-1 ;

  Gij \45:-1 (\P45:31 , \G45:31 , \G30:-1 , \G45:-1 );

  Sum s46(\G45:-1 , A[46], B[46], S[46]);

  wire \P46:45 , \G46:45 ;

  PijGij \46:45 (P[46], P[45], G[46], G[45], \P46:45 , \G46:45 );

  wire \P46:43 , \G46:43 ;

  PijGij \46:43 (\P46:45 , \P44:43 , \G46:45 , \G44:43 , \P46:43 , \G46:43 );

  wire \P46:39 , \G46:39 ;

  PijGij \46:39 (\P46:43 , \P42:39 , \G46:43 , \G42:39 , \P46:39 , \G46:39 );

  wire \P46:31 , \G46:31 ;

  PijGij \46:31 (\P46:39 , \P38:31 , \G46:39 , \G38:31 , \P46:31 , \G46:31 );

  wire \G46:-1 ;

  Gij \46:-1 (\P46:31 , \G46:31 , \G30:-1 , \G46:-1 );

  Sum s47(\G46:-1 , A[47], B[47], S[47]);

  wire \P47:31 , \G47:31 ;

  PijGij \47:31 (P[47], \P46:31 , G[47], \G46:31 , \P47:31 , \G47:31 );

  wire \G47:-1 ;

  Gij \47:-1 (\P47:31 , \G47:31 , \G30:-1 , \G47:-1 );

  Sum s48(\G47:-1 , A[48], B[48], S[48]);

  wire \P48:47 , \G48:47 ;

  PijGij \48:47 (P[48], P[47], G[48], G[47], \P48:47 , \G48:47 );

  wire \P48:31 , \G48:31 ;

  PijGij \48:31 (\P48:47 , \P46:31 , \G48:47 , \G46:31 , \P48:31 , \G48:31 );

  wire \G48:-1 ;

  Gij \48:-1 (\P48:31 , \G48:31 , \G30:-1 , \G48:-1 );

  Sum s49(\G48:-1 , A[49], B[49], S[49]);

  wire \P49:47 , \G49:47 ;

  PijGij \49:47 (P[49], \P48:47 , G[49], \G48:47 , \P49:47 , \G49:47 );

  wire \P49:31 , \G49:31 ;

  PijGij \49:31 (\P49:47 , \P46:31 , \G49:47 , \G46:31 , \P49:31 , \G49:31 );

  wire \G49:-1 ;

  Gij \49:-1 (\P49:31 , \G49:31 , \G30:-1 , \G49:-1 );

  Sum s50(\G49:-1 , A[50], B[50], S[50]);

  wire \P50:49 , \G50:49 ;

  PijGij \50:49 (P[50], P[49], G[50], G[49], \P50:49 , \G50:49 );

  wire \P50:47 , \G50:47 ;

  PijGij \50:47 (\P50:49 , \P48:47 , \G50:49 , \G48:47 , \P50:47 , \G50:47 );

  wire \P50:31 , \G50:31 ;

  PijGij \50:31 (\P50:47 , \P46:31 , \G50:47 , \G46:31 , \P50:31 , \G50:31 );

  wire \G50:-1 ;

  Gij \50:-1 (\P50:31 , \G50:31 , \G30:-1 , \G50:-1 );

  Sum s51(\G50:-1 , A[51], B[51], S[51]);

  wire \P51:47 , \G51:47 ;

  PijGij \51:47 (P[51], \P50:47 , G[51], \G50:47 , \P51:47 , \G51:47 );

  wire \P51:31 , \G51:31 ;

  PijGij \51:31 (\P51:47 , \P46:31 , \G51:47 , \G46:31 , \P51:31 , \G51:31 );

  wire \G51:-1 ;

  Gij \51:-1 (\P51:31 , \G51:31 , \G30:-1 , \G51:-1 );

  Sum s52(\G51:-1 , A[52], B[52], S[52]);

  assign Cout = (\G51:-1 & A[52]) | (\G51:-1 & B[52]) | (A[52] & B[52]);

endmodule
