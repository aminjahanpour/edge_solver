

module padder230(A, B, Cin, S, Cout);
  parameter N = 230;
  input [N-1:0] A, B;
  input Cin;
  output [N-1:0] S;
  output Cout;

  // P[i] is an alias for Pi:i, likewise G[i] is an alias for Gi:i
  wire [N-2:-1] P, G;

  assign P = {A[N-2:0] | B[N-2:0], 1'b0};
  assign G = {A[N-2:0] & B[N-2:0], Cin};

  Sum s0(G[-1], A[0], B[0], S[0]);

  wire \G0:-1 ;

  Gij \0:-1 (P[0], G[0], G[-1], \G0:-1 );

  Sum s1(\G0:-1 , A[1], B[1], S[1]);

  wire \G1:-1 ;

  Gij \1:-1 (P[1], G[1], \G0:-1 , \G1:-1 );

  Sum s2(\G1:-1 , A[2], B[2], S[2]);

  wire \P2:1 , \G2:1 ;

  PijGij \2:1 (P[2], P[1], G[2], G[1], \P2:1 , \G2:1 );

  wire \G2:-1 ;

  Gij \2:-1 (\P2:1 , \G2:1 , \G0:-1 , \G2:-1 );

  Sum s3(\G2:-1 , A[3], B[3], S[3]);

  wire \G3:-1 ;

  Gij \3:-1 (P[3], G[3], \G2:-1 , \G3:-1 );

  Sum s4(\G3:-1 , A[4], B[4], S[4]);

  wire \P4:3 , \G4:3 ;

  PijGij \4:3 (P[4], P[3], G[4], G[3], \P4:3 , \G4:3 );

  wire \G4:-1 ;

  Gij \4:-1 (\P4:3 , \G4:3 , \G2:-1 , \G4:-1 );

  Sum s5(\G4:-1 , A[5], B[5], S[5]);

  wire \P5:3 , \G5:3 ;

  PijGij \5:3 (P[5], \P4:3 , G[5], \G4:3 , \P5:3 , \G5:3 );

  wire \G5:-1 ;

  Gij \5:-1 (\P5:3 , \G5:3 , \G2:-1 , \G5:-1 );

  Sum s6(\G5:-1 , A[6], B[6], S[6]);

  wire \P6:5 , \G6:5 ;

  PijGij \6:5 (P[6], P[5], G[6], G[5], \P6:5 , \G6:5 );

  wire \P6:3 , \G6:3 ;

  PijGij \6:3 (\P6:5 , \P4:3 , \G6:5 , \G4:3 , \P6:3 , \G6:3 );

  wire \G6:-1 ;

  Gij \6:-1 (\P6:3 , \G6:3 , \G2:-1 , \G6:-1 );

  Sum s7(\G6:-1 , A[7], B[7], S[7]);

  wire \G7:-1 ;

  Gij \7:-1 (P[7], G[7], \G6:-1 , \G7:-1 );

  Sum s8(\G7:-1 , A[8], B[8], S[8]);

  wire \P8:7 , \G8:7 ;

  PijGij \8:7 (P[8], P[7], G[8], G[7], \P8:7 , \G8:7 );

  wire \G8:-1 ;

  Gij \8:-1 (\P8:7 , \G8:7 , \G6:-1 , \G8:-1 );

  Sum s9(\G8:-1 , A[9], B[9], S[9]);

  wire \P9:7 , \G9:7 ;

  PijGij \9:7 (P[9], \P8:7 , G[9], \G8:7 , \P9:7 , \G9:7 );

  wire \G9:-1 ;

  Gij \9:-1 (\P9:7 , \G9:7 , \G6:-1 , \G9:-1 );

  Sum s10(\G9:-1 , A[10], B[10], S[10]);

  wire \P10:9 , \G10:9 ;

  PijGij \10:9 (P[10], P[9], G[10], G[9], \P10:9 , \G10:9 );

  wire \P10:7 , \G10:7 ;

  PijGij \10:7 (\P10:9 , \P8:7 , \G10:9 , \G8:7 , \P10:7 , \G10:7 );

  wire \G10:-1 ;

  Gij \10:-1 (\P10:7 , \G10:7 , \G6:-1 , \G10:-1 );

  Sum s11(\G10:-1 , A[11], B[11], S[11]);

  wire \P11:7 , \G11:7 ;

  PijGij \11:7 (P[11], \P10:7 , G[11], \G10:7 , \P11:7 , \G11:7 );

  wire \G11:-1 ;

  Gij \11:-1 (\P11:7 , \G11:7 , \G6:-1 , \G11:-1 );

  Sum s12(\G11:-1 , A[12], B[12], S[12]);

  wire \P12:11 , \G12:11 ;

  PijGij \12:11 (P[12], P[11], G[12], G[11], \P12:11 , \G12:11 );

  wire \P12:7 , \G12:7 ;

  PijGij \12:7 (\P12:11 , \P10:7 , \G12:11 , \G10:7 , \P12:7 , \G12:7 );

  wire \G12:-1 ;

  Gij \12:-1 (\P12:7 , \G12:7 , \G6:-1 , \G12:-1 );

  Sum s13(\G12:-1 , A[13], B[13], S[13]);

  wire \P13:11 , \G13:11 ;

  PijGij \13:11 (P[13], \P12:11 , G[13], \G12:11 , \P13:11 , \G13:11 );

  wire \P13:7 , \G13:7 ;

  PijGij \13:7 (\P13:11 , \P10:7 , \G13:11 , \G10:7 , \P13:7 , \G13:7 );

  wire \G13:-1 ;

  Gij \13:-1 (\P13:7 , \G13:7 , \G6:-1 , \G13:-1 );

  Sum s14(\G13:-1 , A[14], B[14], S[14]);

  wire \P14:13 , \G14:13 ;

  PijGij \14:13 (P[14], P[13], G[14], G[13], \P14:13 , \G14:13 );

  wire \P14:11 , \G14:11 ;

  PijGij \14:11 (\P14:13 , \P12:11 , \G14:13 , \G12:11 , \P14:11 , \G14:11 );

  wire \P14:7 , \G14:7 ;

  PijGij \14:7 (\P14:11 , \P10:7 , \G14:11 , \G10:7 , \P14:7 , \G14:7 );

  wire \G14:-1 ;

  Gij \14:-1 (\P14:7 , \G14:7 , \G6:-1 , \G14:-1 );

  Sum s15(\G14:-1 , A[15], B[15], S[15]);

  wire \G15:-1 ;

  Gij \15:-1 (P[15], G[15], \G14:-1 , \G15:-1 );

  Sum s16(\G15:-1 , A[16], B[16], S[16]);

  wire \P16:15 , \G16:15 ;

  PijGij \16:15 (P[16], P[15], G[16], G[15], \P16:15 , \G16:15 );

  wire \G16:-1 ;

  Gij \16:-1 (\P16:15 , \G16:15 , \G14:-1 , \G16:-1 );

  Sum s17(\G16:-1 , A[17], B[17], S[17]);

  wire \P17:15 , \G17:15 ;

  PijGij \17:15 (P[17], \P16:15 , G[17], \G16:15 , \P17:15 , \G17:15 );

  wire \G17:-1 ;

  Gij \17:-1 (\P17:15 , \G17:15 , \G14:-1 , \G17:-1 );

  Sum s18(\G17:-1 , A[18], B[18], S[18]);

  wire \P18:17 , \G18:17 ;

  PijGij \18:17 (P[18], P[17], G[18], G[17], \P18:17 , \G18:17 );

  wire \P18:15 , \G18:15 ;

  PijGij \18:15 (\P18:17 , \P16:15 , \G18:17 , \G16:15 , \P18:15 , \G18:15 );

  wire \G18:-1 ;

  Gij \18:-1 (\P18:15 , \G18:15 , \G14:-1 , \G18:-1 );

  Sum s19(\G18:-1 , A[19], B[19], S[19]);

  wire \P19:15 , \G19:15 ;

  PijGij \19:15 (P[19], \P18:15 , G[19], \G18:15 , \P19:15 , \G19:15 );

  wire \G19:-1 ;

  Gij \19:-1 (\P19:15 , \G19:15 , \G14:-1 , \G19:-1 );

  Sum s20(\G19:-1 , A[20], B[20], S[20]);

  wire \P20:19 , \G20:19 ;

  PijGij \20:19 (P[20], P[19], G[20], G[19], \P20:19 , \G20:19 );

  wire \P20:15 , \G20:15 ;

  PijGij \20:15 (\P20:19 , \P18:15 , \G20:19 , \G18:15 , \P20:15 , \G20:15 );

  wire \G20:-1 ;

  Gij \20:-1 (\P20:15 , \G20:15 , \G14:-1 , \G20:-1 );

  Sum s21(\G20:-1 , A[21], B[21], S[21]);

  wire \P21:19 , \G21:19 ;

  PijGij \21:19 (P[21], \P20:19 , G[21], \G20:19 , \P21:19 , \G21:19 );

  wire \P21:15 , \G21:15 ;

  PijGij \21:15 (\P21:19 , \P18:15 , \G21:19 , \G18:15 , \P21:15 , \G21:15 );

  wire \G21:-1 ;

  Gij \21:-1 (\P21:15 , \G21:15 , \G14:-1 , \G21:-1 );

  Sum s22(\G21:-1 , A[22], B[22], S[22]);

  wire \P22:21 , \G22:21 ;

  PijGij \22:21 (P[22], P[21], G[22], G[21], \P22:21 , \G22:21 );

  wire \P22:19 , \G22:19 ;

  PijGij \22:19 (\P22:21 , \P20:19 , \G22:21 , \G20:19 , \P22:19 , \G22:19 );

  wire \P22:15 , \G22:15 ;

  PijGij \22:15 (\P22:19 , \P18:15 , \G22:19 , \G18:15 , \P22:15 , \G22:15 );

  wire \G22:-1 ;

  Gij \22:-1 (\P22:15 , \G22:15 , \G14:-1 , \G22:-1 );

  Sum s23(\G22:-1 , A[23], B[23], S[23]);

  wire \P23:15 , \G23:15 ;

  PijGij \23:15 (P[23], \P22:15 , G[23], \G22:15 , \P23:15 , \G23:15 );

  wire \G23:-1 ;

  Gij \23:-1 (\P23:15 , \G23:15 , \G14:-1 , \G23:-1 );

  Sum s24(\G23:-1 , A[24], B[24], S[24]);

  wire \P24:23 , \G24:23 ;

  PijGij \24:23 (P[24], P[23], G[24], G[23], \P24:23 , \G24:23 );

  wire \P24:15 , \G24:15 ;

  PijGij \24:15 (\P24:23 , \P22:15 , \G24:23 , \G22:15 , \P24:15 , \G24:15 );

  wire \G24:-1 ;

  Gij \24:-1 (\P24:15 , \G24:15 , \G14:-1 , \G24:-1 );

  Sum s25(\G24:-1 , A[25], B[25], S[25]);

  wire \P25:23 , \G25:23 ;

  PijGij \25:23 (P[25], \P24:23 , G[25], \G24:23 , \P25:23 , \G25:23 );

  wire \P25:15 , \G25:15 ;

  PijGij \25:15 (\P25:23 , \P22:15 , \G25:23 , \G22:15 , \P25:15 , \G25:15 );

  wire \G25:-1 ;

  Gij \25:-1 (\P25:15 , \G25:15 , \G14:-1 , \G25:-1 );

  Sum s26(\G25:-1 , A[26], B[26], S[26]);

  wire \P26:25 , \G26:25 ;

  PijGij \26:25 (P[26], P[25], G[26], G[25], \P26:25 , \G26:25 );

  wire \P26:23 , \G26:23 ;

  PijGij \26:23 (\P26:25 , \P24:23 , \G26:25 , \G24:23 , \P26:23 , \G26:23 );

  wire \P26:15 , \G26:15 ;

  PijGij \26:15 (\P26:23 , \P22:15 , \G26:23 , \G22:15 , \P26:15 , \G26:15 );

  wire \G26:-1 ;

  Gij \26:-1 (\P26:15 , \G26:15 , \G14:-1 , \G26:-1 );

  Sum s27(\G26:-1 , A[27], B[27], S[27]);

  wire \P27:23 , \G27:23 ;

  PijGij \27:23 (P[27], \P26:23 , G[27], \G26:23 , \P27:23 , \G27:23 );

  wire \P27:15 , \G27:15 ;

  PijGij \27:15 (\P27:23 , \P22:15 , \G27:23 , \G22:15 , \P27:15 , \G27:15 );

  wire \G27:-1 ;

  Gij \27:-1 (\P27:15 , \G27:15 , \G14:-1 , \G27:-1 );

  Sum s28(\G27:-1 , A[28], B[28], S[28]);

  wire \P28:27 , \G28:27 ;

  PijGij \28:27 (P[28], P[27], G[28], G[27], \P28:27 , \G28:27 );

  wire \P28:23 , \G28:23 ;

  PijGij \28:23 (\P28:27 , \P26:23 , \G28:27 , \G26:23 , \P28:23 , \G28:23 );

  wire \P28:15 , \G28:15 ;

  PijGij \28:15 (\P28:23 , \P22:15 , \G28:23 , \G22:15 , \P28:15 , \G28:15 );

  wire \G28:-1 ;

  Gij \28:-1 (\P28:15 , \G28:15 , \G14:-1 , \G28:-1 );

  Sum s29(\G28:-1 , A[29], B[29], S[29]);

  wire \P29:27 , \G29:27 ;

  PijGij \29:27 (P[29], \P28:27 , G[29], \G28:27 , \P29:27 , \G29:27 );

  wire \P29:23 , \G29:23 ;

  PijGij \29:23 (\P29:27 , \P26:23 , \G29:27 , \G26:23 , \P29:23 , \G29:23 );

  wire \P29:15 , \G29:15 ;

  PijGij \29:15 (\P29:23 , \P22:15 , \G29:23 , \G22:15 , \P29:15 , \G29:15 );

  wire \G29:-1 ;

  Gij \29:-1 (\P29:15 , \G29:15 , \G14:-1 , \G29:-1 );

  Sum s30(\G29:-1 , A[30], B[30], S[30]);

  wire \P30:29 , \G30:29 ;

  PijGij \30:29 (P[30], P[29], G[30], G[29], \P30:29 , \G30:29 );

  wire \P30:27 , \G30:27 ;

  PijGij \30:27 (\P30:29 , \P28:27 , \G30:29 , \G28:27 , \P30:27 , \G30:27 );

  wire \P30:23 , \G30:23 ;

  PijGij \30:23 (\P30:27 , \P26:23 , \G30:27 , \G26:23 , \P30:23 , \G30:23 );

  wire \P30:15 , \G30:15 ;

  PijGij \30:15 (\P30:23 , \P22:15 , \G30:23 , \G22:15 , \P30:15 , \G30:15 );

  wire \G30:-1 ;

  Gij \30:-1 (\P30:15 , \G30:15 , \G14:-1 , \G30:-1 );

  Sum s31(\G30:-1 , A[31], B[31], S[31]);

  wire \G31:-1 ;

  Gij \31:-1 (P[31], G[31], \G30:-1 , \G31:-1 );

  Sum s32(\G31:-1 , A[32], B[32], S[32]);

  wire \P32:31 , \G32:31 ;

  PijGij \32:31 (P[32], P[31], G[32], G[31], \P32:31 , \G32:31 );

  wire \G32:-1 ;

  Gij \32:-1 (\P32:31 , \G32:31 , \G30:-1 , \G32:-1 );

  Sum s33(\G32:-1 , A[33], B[33], S[33]);

  wire \P33:31 , \G33:31 ;

  PijGij \33:31 (P[33], \P32:31 , G[33], \G32:31 , \P33:31 , \G33:31 );

  wire \G33:-1 ;

  Gij \33:-1 (\P33:31 , \G33:31 , \G30:-1 , \G33:-1 );

  Sum s34(\G33:-1 , A[34], B[34], S[34]);

  wire \P34:33 , \G34:33 ;

  PijGij \34:33 (P[34], P[33], G[34], G[33], \P34:33 , \G34:33 );

  wire \P34:31 , \G34:31 ;

  PijGij \34:31 (\P34:33 , \P32:31 , \G34:33 , \G32:31 , \P34:31 , \G34:31 );

  wire \G34:-1 ;

  Gij \34:-1 (\P34:31 , \G34:31 , \G30:-1 , \G34:-1 );

  Sum s35(\G34:-1 , A[35], B[35], S[35]);

  wire \P35:31 , \G35:31 ;

  PijGij \35:31 (P[35], \P34:31 , G[35], \G34:31 , \P35:31 , \G35:31 );

  wire \G35:-1 ;

  Gij \35:-1 (\P35:31 , \G35:31 , \G30:-1 , \G35:-1 );

  Sum s36(\G35:-1 , A[36], B[36], S[36]);

  wire \P36:35 , \G36:35 ;

  PijGij \36:35 (P[36], P[35], G[36], G[35], \P36:35 , \G36:35 );

  wire \P36:31 , \G36:31 ;

  PijGij \36:31 (\P36:35 , \P34:31 , \G36:35 , \G34:31 , \P36:31 , \G36:31 );

  wire \G36:-1 ;

  Gij \36:-1 (\P36:31 , \G36:31 , \G30:-1 , \G36:-1 );

  Sum s37(\G36:-1 , A[37], B[37], S[37]);

  wire \P37:35 , \G37:35 ;

  PijGij \37:35 (P[37], \P36:35 , G[37], \G36:35 , \P37:35 , \G37:35 );

  wire \P37:31 , \G37:31 ;

  PijGij \37:31 (\P37:35 , \P34:31 , \G37:35 , \G34:31 , \P37:31 , \G37:31 );

  wire \G37:-1 ;

  Gij \37:-1 (\P37:31 , \G37:31 , \G30:-1 , \G37:-1 );

  Sum s38(\G37:-1 , A[38], B[38], S[38]);

  wire \P38:37 , \G38:37 ;

  PijGij \38:37 (P[38], P[37], G[38], G[37], \P38:37 , \G38:37 );

  wire \P38:35 , \G38:35 ;

  PijGij \38:35 (\P38:37 , \P36:35 , \G38:37 , \G36:35 , \P38:35 , \G38:35 );

  wire \P38:31 , \G38:31 ;

  PijGij \38:31 (\P38:35 , \P34:31 , \G38:35 , \G34:31 , \P38:31 , \G38:31 );

  wire \G38:-1 ;

  Gij \38:-1 (\P38:31 , \G38:31 , \G30:-1 , \G38:-1 );

  Sum s39(\G38:-1 , A[39], B[39], S[39]);

  wire \P39:31 , \G39:31 ;

  PijGij \39:31 (P[39], \P38:31 , G[39], \G38:31 , \P39:31 , \G39:31 );

  wire \G39:-1 ;

  Gij \39:-1 (\P39:31 , \G39:31 , \G30:-1 , \G39:-1 );

  Sum s40(\G39:-1 , A[40], B[40], S[40]);

  wire \P40:39 , \G40:39 ;

  PijGij \40:39 (P[40], P[39], G[40], G[39], \P40:39 , \G40:39 );

  wire \P40:31 , \G40:31 ;

  PijGij \40:31 (\P40:39 , \P38:31 , \G40:39 , \G38:31 , \P40:31 , \G40:31 );

  wire \G40:-1 ;

  Gij \40:-1 (\P40:31 , \G40:31 , \G30:-1 , \G40:-1 );

  Sum s41(\G40:-1 , A[41], B[41], S[41]);

  wire \P41:39 , \G41:39 ;

  PijGij \41:39 (P[41], \P40:39 , G[41], \G40:39 , \P41:39 , \G41:39 );

  wire \P41:31 , \G41:31 ;

  PijGij \41:31 (\P41:39 , \P38:31 , \G41:39 , \G38:31 , \P41:31 , \G41:31 );

  wire \G41:-1 ;

  Gij \41:-1 (\P41:31 , \G41:31 , \G30:-1 , \G41:-1 );

  Sum s42(\G41:-1 , A[42], B[42], S[42]);

  wire \P42:41 , \G42:41 ;

  PijGij \42:41 (P[42], P[41], G[42], G[41], \P42:41 , \G42:41 );

  wire \P42:39 , \G42:39 ;

  PijGij \42:39 (\P42:41 , \P40:39 , \G42:41 , \G40:39 , \P42:39 , \G42:39 );

  wire \P42:31 , \G42:31 ;

  PijGij \42:31 (\P42:39 , \P38:31 , \G42:39 , \G38:31 , \P42:31 , \G42:31 );

  wire \G42:-1 ;

  Gij \42:-1 (\P42:31 , \G42:31 , \G30:-1 , \G42:-1 );

  Sum s43(\G42:-1 , A[43], B[43], S[43]);

  wire \P43:39 , \G43:39 ;

  PijGij \43:39 (P[43], \P42:39 , G[43], \G42:39 , \P43:39 , \G43:39 );

  wire \P43:31 , \G43:31 ;

  PijGij \43:31 (\P43:39 , \P38:31 , \G43:39 , \G38:31 , \P43:31 , \G43:31 );

  wire \G43:-1 ;

  Gij \43:-1 (\P43:31 , \G43:31 , \G30:-1 , \G43:-1 );

  Sum s44(\G43:-1 , A[44], B[44], S[44]);

  wire \P44:43 , \G44:43 ;

  PijGij \44:43 (P[44], P[43], G[44], G[43], \P44:43 , \G44:43 );

  wire \P44:39 , \G44:39 ;

  PijGij \44:39 (\P44:43 , \P42:39 , \G44:43 , \G42:39 , \P44:39 , \G44:39 );

  wire \P44:31 , \G44:31 ;

  PijGij \44:31 (\P44:39 , \P38:31 , \G44:39 , \G38:31 , \P44:31 , \G44:31 );

  wire \G44:-1 ;

  Gij \44:-1 (\P44:31 , \G44:31 , \G30:-1 , \G44:-1 );

  Sum s45(\G44:-1 , A[45], B[45], S[45]);

  wire \P45:43 , \G45:43 ;

  PijGij \45:43 (P[45], \P44:43 , G[45], \G44:43 , \P45:43 , \G45:43 );

  wire \P45:39 , \G45:39 ;

  PijGij \45:39 (\P45:43 , \P42:39 , \G45:43 , \G42:39 , \P45:39 , \G45:39 );

  wire \P45:31 , \G45:31 ;

  PijGij \45:31 (\P45:39 , \P38:31 , \G45:39 , \G38:31 , \P45:31 , \G45:31 );

  wire \G45:-1 ;

  Gij \45:-1 (\P45:31 , \G45:31 , \G30:-1 , \G45:-1 );

  Sum s46(\G45:-1 , A[46], B[46], S[46]);

  wire \P46:45 , \G46:45 ;

  PijGij \46:45 (P[46], P[45], G[46], G[45], \P46:45 , \G46:45 );

  wire \P46:43 , \G46:43 ;

  PijGij \46:43 (\P46:45 , \P44:43 , \G46:45 , \G44:43 , \P46:43 , \G46:43 );

  wire \P46:39 , \G46:39 ;

  PijGij \46:39 (\P46:43 , \P42:39 , \G46:43 , \G42:39 , \P46:39 , \G46:39 );

  wire \P46:31 , \G46:31 ;

  PijGij \46:31 (\P46:39 , \P38:31 , \G46:39 , \G38:31 , \P46:31 , \G46:31 );

  wire \G46:-1 ;

  Gij \46:-1 (\P46:31 , \G46:31 , \G30:-1 , \G46:-1 );

  Sum s47(\G46:-1 , A[47], B[47], S[47]);

  wire \P47:31 , \G47:31 ;

  PijGij \47:31 (P[47], \P46:31 , G[47], \G46:31 , \P47:31 , \G47:31 );

  wire \G47:-1 ;

  Gij \47:-1 (\P47:31 , \G47:31 , \G30:-1 , \G47:-1 );

  Sum s48(\G47:-1 , A[48], B[48], S[48]);

  wire \P48:47 , \G48:47 ;

  PijGij \48:47 (P[48], P[47], G[48], G[47], \P48:47 , \G48:47 );

  wire \P48:31 , \G48:31 ;

  PijGij \48:31 (\P48:47 , \P46:31 , \G48:47 , \G46:31 , \P48:31 , \G48:31 );

  wire \G48:-1 ;

  Gij \48:-1 (\P48:31 , \G48:31 , \G30:-1 , \G48:-1 );

  Sum s49(\G48:-1 , A[49], B[49], S[49]);

  wire \P49:47 , \G49:47 ;

  PijGij \49:47 (P[49], \P48:47 , G[49], \G48:47 , \P49:47 , \G49:47 );

  wire \P49:31 , \G49:31 ;

  PijGij \49:31 (\P49:47 , \P46:31 , \G49:47 , \G46:31 , \P49:31 , \G49:31 );

  wire \G49:-1 ;

  Gij \49:-1 (\P49:31 , \G49:31 , \G30:-1 , \G49:-1 );

  Sum s50(\G49:-1 , A[50], B[50], S[50]);

  wire \P50:49 , \G50:49 ;

  PijGij \50:49 (P[50], P[49], G[50], G[49], \P50:49 , \G50:49 );

  wire \P50:47 , \G50:47 ;

  PijGij \50:47 (\P50:49 , \P48:47 , \G50:49 , \G48:47 , \P50:47 , \G50:47 );

  wire \P50:31 , \G50:31 ;

  PijGij \50:31 (\P50:47 , \P46:31 , \G50:47 , \G46:31 , \P50:31 , \G50:31 );

  wire \G50:-1 ;

  Gij \50:-1 (\P50:31 , \G50:31 , \G30:-1 , \G50:-1 );

  Sum s51(\G50:-1 , A[51], B[51], S[51]);

  wire \P51:47 , \G51:47 ;

  PijGij \51:47 (P[51], \P50:47 , G[51], \G50:47 , \P51:47 , \G51:47 );

  wire \P51:31 , \G51:31 ;

  PijGij \51:31 (\P51:47 , \P46:31 , \G51:47 , \G46:31 , \P51:31 , \G51:31 );

  wire \G51:-1 ;

  Gij \51:-1 (\P51:31 , \G51:31 , \G30:-1 , \G51:-1 );

  Sum s52(\G51:-1 , A[52], B[52], S[52]);

  wire \P52:51 , \G52:51 ;

  PijGij \52:51 (P[52], P[51], G[52], G[51], \P52:51 , \G52:51 );

  wire \P52:47 , \G52:47 ;

  PijGij \52:47 (\P52:51 , \P50:47 , \G52:51 , \G50:47 , \P52:47 , \G52:47 );

  wire \P52:31 , \G52:31 ;

  PijGij \52:31 (\P52:47 , \P46:31 , \G52:47 , \G46:31 , \P52:31 , \G52:31 );

  wire \G52:-1 ;

  Gij \52:-1 (\P52:31 , \G52:31 , \G30:-1 , \G52:-1 );

  Sum s53(\G52:-1 , A[53], B[53], S[53]);

  wire \P53:51 , \G53:51 ;

  PijGij \53:51 (P[53], \P52:51 , G[53], \G52:51 , \P53:51 , \G53:51 );

  wire \P53:47 , \G53:47 ;

  PijGij \53:47 (\P53:51 , \P50:47 , \G53:51 , \G50:47 , \P53:47 , \G53:47 );

  wire \P53:31 , \G53:31 ;

  PijGij \53:31 (\P53:47 , \P46:31 , \G53:47 , \G46:31 , \P53:31 , \G53:31 );

  wire \G53:-1 ;

  Gij \53:-1 (\P53:31 , \G53:31 , \G30:-1 , \G53:-1 );

  Sum s54(\G53:-1 , A[54], B[54], S[54]);

  wire \P54:53 , \G54:53 ;

  PijGij \54:53 (P[54], P[53], G[54], G[53], \P54:53 , \G54:53 );

  wire \P54:51 , \G54:51 ;

  PijGij \54:51 (\P54:53 , \P52:51 , \G54:53 , \G52:51 , \P54:51 , \G54:51 );

  wire \P54:47 , \G54:47 ;

  PijGij \54:47 (\P54:51 , \P50:47 , \G54:51 , \G50:47 , \P54:47 , \G54:47 );

  wire \P54:31 , \G54:31 ;

  PijGij \54:31 (\P54:47 , \P46:31 , \G54:47 , \G46:31 , \P54:31 , \G54:31 );

  wire \G54:-1 ;

  Gij \54:-1 (\P54:31 , \G54:31 , \G30:-1 , \G54:-1 );

  Sum s55(\G54:-1 , A[55], B[55], S[55]);

  wire \P55:47 , \G55:47 ;

  PijGij \55:47 (P[55], \P54:47 , G[55], \G54:47 , \P55:47 , \G55:47 );

  wire \P55:31 , \G55:31 ;

  PijGij \55:31 (\P55:47 , \P46:31 , \G55:47 , \G46:31 , \P55:31 , \G55:31 );

  wire \G55:-1 ;

  Gij \55:-1 (\P55:31 , \G55:31 , \G30:-1 , \G55:-1 );

  Sum s56(\G55:-1 , A[56], B[56], S[56]);

  wire \P56:55 , \G56:55 ;

  PijGij \56:55 (P[56], P[55], G[56], G[55], \P56:55 , \G56:55 );

  wire \P56:47 , \G56:47 ;

  PijGij \56:47 (\P56:55 , \P54:47 , \G56:55 , \G54:47 , \P56:47 , \G56:47 );

  wire \P56:31 , \G56:31 ;

  PijGij \56:31 (\P56:47 , \P46:31 , \G56:47 , \G46:31 , \P56:31 , \G56:31 );

  wire \G56:-1 ;

  Gij \56:-1 (\P56:31 , \G56:31 , \G30:-1 , \G56:-1 );

  Sum s57(\G56:-1 , A[57], B[57], S[57]);

  wire \P57:55 , \G57:55 ;

  PijGij \57:55 (P[57], \P56:55 , G[57], \G56:55 , \P57:55 , \G57:55 );

  wire \P57:47 , \G57:47 ;

  PijGij \57:47 (\P57:55 , \P54:47 , \G57:55 , \G54:47 , \P57:47 , \G57:47 );

  wire \P57:31 , \G57:31 ;

  PijGij \57:31 (\P57:47 , \P46:31 , \G57:47 , \G46:31 , \P57:31 , \G57:31 );

  wire \G57:-1 ;

  Gij \57:-1 (\P57:31 , \G57:31 , \G30:-1 , \G57:-1 );

  Sum s58(\G57:-1 , A[58], B[58], S[58]);

  wire \P58:57 , \G58:57 ;

  PijGij \58:57 (P[58], P[57], G[58], G[57], \P58:57 , \G58:57 );

  wire \P58:55 , \G58:55 ;

  PijGij \58:55 (\P58:57 , \P56:55 , \G58:57 , \G56:55 , \P58:55 , \G58:55 );

  wire \P58:47 , \G58:47 ;

  PijGij \58:47 (\P58:55 , \P54:47 , \G58:55 , \G54:47 , \P58:47 , \G58:47 );

  wire \P58:31 , \G58:31 ;

  PijGij \58:31 (\P58:47 , \P46:31 , \G58:47 , \G46:31 , \P58:31 , \G58:31 );

  wire \G58:-1 ;

  Gij \58:-1 (\P58:31 , \G58:31 , \G30:-1 , \G58:-1 );

  Sum s59(\G58:-1 , A[59], B[59], S[59]);

  wire \P59:55 , \G59:55 ;

  PijGij \59:55 (P[59], \P58:55 , G[59], \G58:55 , \P59:55 , \G59:55 );

  wire \P59:47 , \G59:47 ;

  PijGij \59:47 (\P59:55 , \P54:47 , \G59:55 , \G54:47 , \P59:47 , \G59:47 );

  wire \P59:31 , \G59:31 ;

  PijGij \59:31 (\P59:47 , \P46:31 , \G59:47 , \G46:31 , \P59:31 , \G59:31 );

  wire \G59:-1 ;

  Gij \59:-1 (\P59:31 , \G59:31 , \G30:-1 , \G59:-1 );

  Sum s60(\G59:-1 , A[60], B[60], S[60]);

  wire \P60:59 , \G60:59 ;

  PijGij \60:59 (P[60], P[59], G[60], G[59], \P60:59 , \G60:59 );

  wire \P60:55 , \G60:55 ;

  PijGij \60:55 (\P60:59 , \P58:55 , \G60:59 , \G58:55 , \P60:55 , \G60:55 );

  wire \P60:47 , \G60:47 ;

  PijGij \60:47 (\P60:55 , \P54:47 , \G60:55 , \G54:47 , \P60:47 , \G60:47 );

  wire \P60:31 , \G60:31 ;

  PijGij \60:31 (\P60:47 , \P46:31 , \G60:47 , \G46:31 , \P60:31 , \G60:31 );

  wire \G60:-1 ;

  Gij \60:-1 (\P60:31 , \G60:31 , \G30:-1 , \G60:-1 );

  Sum s61(\G60:-1 , A[61], B[61], S[61]);

  wire \P61:59 , \G61:59 ;

  PijGij \61:59 (P[61], \P60:59 , G[61], \G60:59 , \P61:59 , \G61:59 );

  wire \P61:55 , \G61:55 ;

  PijGij \61:55 (\P61:59 , \P58:55 , \G61:59 , \G58:55 , \P61:55 , \G61:55 );

  wire \P61:47 , \G61:47 ;

  PijGij \61:47 (\P61:55 , \P54:47 , \G61:55 , \G54:47 , \P61:47 , \G61:47 );

  wire \P61:31 , \G61:31 ;

  PijGij \61:31 (\P61:47 , \P46:31 , \G61:47 , \G46:31 , \P61:31 , \G61:31 );

  wire \G61:-1 ;

  Gij \61:-1 (\P61:31 , \G61:31 , \G30:-1 , \G61:-1 );

  Sum s62(\G61:-1 , A[62], B[62], S[62]);

  wire \P62:61 , \G62:61 ;

  PijGij \62:61 (P[62], P[61], G[62], G[61], \P62:61 , \G62:61 );

  wire \P62:59 , \G62:59 ;

  PijGij \62:59 (\P62:61 , \P60:59 , \G62:61 , \G60:59 , \P62:59 , \G62:59 );

  wire \P62:55 , \G62:55 ;

  PijGij \62:55 (\P62:59 , \P58:55 , \G62:59 , \G58:55 , \P62:55 , \G62:55 );

  wire \P62:47 , \G62:47 ;

  PijGij \62:47 (\P62:55 , \P54:47 , \G62:55 , \G54:47 , \P62:47 , \G62:47 );

  wire \P62:31 , \G62:31 ;

  PijGij \62:31 (\P62:47 , \P46:31 , \G62:47 , \G46:31 , \P62:31 , \G62:31 );

  wire \G62:-1 ;

  Gij \62:-1 (\P62:31 , \G62:31 , \G30:-1 , \G62:-1 );

  Sum s63(\G62:-1 , A[63], B[63], S[63]);

  wire \G63:-1 ;

  Gij \63:-1 (P[63], G[63], \G62:-1 , \G63:-1 );

  Sum s64(\G63:-1 , A[64], B[64], S[64]);

  wire \P64:63 , \G64:63 ;

  PijGij \64:63 (P[64], P[63], G[64], G[63], \P64:63 , \G64:63 );

  wire \G64:-1 ;

  Gij \64:-1 (\P64:63 , \G64:63 , \G62:-1 , \G64:-1 );

  Sum s65(\G64:-1 , A[65], B[65], S[65]);

  wire \P65:63 , \G65:63 ;

  PijGij \65:63 (P[65], \P64:63 , G[65], \G64:63 , \P65:63 , \G65:63 );

  wire \G65:-1 ;

  Gij \65:-1 (\P65:63 , \G65:63 , \G62:-1 , \G65:-1 );

  Sum s66(\G65:-1 , A[66], B[66], S[66]);

  wire \P66:65 , \G66:65 ;

  PijGij \66:65 (P[66], P[65], G[66], G[65], \P66:65 , \G66:65 );

  wire \P66:63 , \G66:63 ;

  PijGij \66:63 (\P66:65 , \P64:63 , \G66:65 , \G64:63 , \P66:63 , \G66:63 );

  wire \G66:-1 ;

  Gij \66:-1 (\P66:63 , \G66:63 , \G62:-1 , \G66:-1 );

  Sum s67(\G66:-1 , A[67], B[67], S[67]);

  wire \P67:63 , \G67:63 ;

  PijGij \67:63 (P[67], \P66:63 , G[67], \G66:63 , \P67:63 , \G67:63 );

  wire \G67:-1 ;

  Gij \67:-1 (\P67:63 , \G67:63 , \G62:-1 , \G67:-1 );

  Sum s68(\G67:-1 , A[68], B[68], S[68]);

  wire \P68:67 , \G68:67 ;

  PijGij \68:67 (P[68], P[67], G[68], G[67], \P68:67 , \G68:67 );

  wire \P68:63 , \G68:63 ;

  PijGij \68:63 (\P68:67 , \P66:63 , \G68:67 , \G66:63 , \P68:63 , \G68:63 );

  wire \G68:-1 ;

  Gij \68:-1 (\P68:63 , \G68:63 , \G62:-1 , \G68:-1 );

  Sum s69(\G68:-1 , A[69], B[69], S[69]);

  wire \P69:67 , \G69:67 ;

  PijGij \69:67 (P[69], \P68:67 , G[69], \G68:67 , \P69:67 , \G69:67 );

  wire \P69:63 , \G69:63 ;

  PijGij \69:63 (\P69:67 , \P66:63 , \G69:67 , \G66:63 , \P69:63 , \G69:63 );

  wire \G69:-1 ;

  Gij \69:-1 (\P69:63 , \G69:63 , \G62:-1 , \G69:-1 );

  Sum s70(\G69:-1 , A[70], B[70], S[70]);

  wire \P70:69 , \G70:69 ;

  PijGij \70:69 (P[70], P[69], G[70], G[69], \P70:69 , \G70:69 );

  wire \P70:67 , \G70:67 ;

  PijGij \70:67 (\P70:69 , \P68:67 , \G70:69 , \G68:67 , \P70:67 , \G70:67 );

  wire \P70:63 , \G70:63 ;

  PijGij \70:63 (\P70:67 , \P66:63 , \G70:67 , \G66:63 , \P70:63 , \G70:63 );

  wire \G70:-1 ;

  Gij \70:-1 (\P70:63 , \G70:63 , \G62:-1 , \G70:-1 );

  Sum s71(\G70:-1 , A[71], B[71], S[71]);

  wire \P71:63 , \G71:63 ;

  PijGij \71:63 (P[71], \P70:63 , G[71], \G70:63 , \P71:63 , \G71:63 );

  wire \G71:-1 ;

  Gij \71:-1 (\P71:63 , \G71:63 , \G62:-1 , \G71:-1 );

  Sum s72(\G71:-1 , A[72], B[72], S[72]);

  wire \P72:71 , \G72:71 ;

  PijGij \72:71 (P[72], P[71], G[72], G[71], \P72:71 , \G72:71 );

  wire \P72:63 , \G72:63 ;

  PijGij \72:63 (\P72:71 , \P70:63 , \G72:71 , \G70:63 , \P72:63 , \G72:63 );

  wire \G72:-1 ;

  Gij \72:-1 (\P72:63 , \G72:63 , \G62:-1 , \G72:-1 );

  Sum s73(\G72:-1 , A[73], B[73], S[73]);

  wire \P73:71 , \G73:71 ;

  PijGij \73:71 (P[73], \P72:71 , G[73], \G72:71 , \P73:71 , \G73:71 );

  wire \P73:63 , \G73:63 ;

  PijGij \73:63 (\P73:71 , \P70:63 , \G73:71 , \G70:63 , \P73:63 , \G73:63 );

  wire \G73:-1 ;

  Gij \73:-1 (\P73:63 , \G73:63 , \G62:-1 , \G73:-1 );

  Sum s74(\G73:-1 , A[74], B[74], S[74]);

  wire \P74:73 , \G74:73 ;

  PijGij \74:73 (P[74], P[73], G[74], G[73], \P74:73 , \G74:73 );

  wire \P74:71 , \G74:71 ;

  PijGij \74:71 (\P74:73 , \P72:71 , \G74:73 , \G72:71 , \P74:71 , \G74:71 );

  wire \P74:63 , \G74:63 ;

  PijGij \74:63 (\P74:71 , \P70:63 , \G74:71 , \G70:63 , \P74:63 , \G74:63 );

  wire \G74:-1 ;

  Gij \74:-1 (\P74:63 , \G74:63 , \G62:-1 , \G74:-1 );

  Sum s75(\G74:-1 , A[75], B[75], S[75]);

  wire \P75:71 , \G75:71 ;

  PijGij \75:71 (P[75], \P74:71 , G[75], \G74:71 , \P75:71 , \G75:71 );

  wire \P75:63 , \G75:63 ;

  PijGij \75:63 (\P75:71 , \P70:63 , \G75:71 , \G70:63 , \P75:63 , \G75:63 );

  wire \G75:-1 ;

  Gij \75:-1 (\P75:63 , \G75:63 , \G62:-1 , \G75:-1 );

  Sum s76(\G75:-1 , A[76], B[76], S[76]);

  wire \P76:75 , \G76:75 ;

  PijGij \76:75 (P[76], P[75], G[76], G[75], \P76:75 , \G76:75 );

  wire \P76:71 , \G76:71 ;

  PijGij \76:71 (\P76:75 , \P74:71 , \G76:75 , \G74:71 , \P76:71 , \G76:71 );

  wire \P76:63 , \G76:63 ;

  PijGij \76:63 (\P76:71 , \P70:63 , \G76:71 , \G70:63 , \P76:63 , \G76:63 );

  wire \G76:-1 ;

  Gij \76:-1 (\P76:63 , \G76:63 , \G62:-1 , \G76:-1 );

  Sum s77(\G76:-1 , A[77], B[77], S[77]);

  wire \P77:75 , \G77:75 ;

  PijGij \77:75 (P[77], \P76:75 , G[77], \G76:75 , \P77:75 , \G77:75 );

  wire \P77:71 , \G77:71 ;

  PijGij \77:71 (\P77:75 , \P74:71 , \G77:75 , \G74:71 , \P77:71 , \G77:71 );

  wire \P77:63 , \G77:63 ;

  PijGij \77:63 (\P77:71 , \P70:63 , \G77:71 , \G70:63 , \P77:63 , \G77:63 );

  wire \G77:-1 ;

  Gij \77:-1 (\P77:63 , \G77:63 , \G62:-1 , \G77:-1 );

  Sum s78(\G77:-1 , A[78], B[78], S[78]);

  wire \P78:77 , \G78:77 ;

  PijGij \78:77 (P[78], P[77], G[78], G[77], \P78:77 , \G78:77 );

  wire \P78:75 , \G78:75 ;

  PijGij \78:75 (\P78:77 , \P76:75 , \G78:77 , \G76:75 , \P78:75 , \G78:75 );

  wire \P78:71 , \G78:71 ;

  PijGij \78:71 (\P78:75 , \P74:71 , \G78:75 , \G74:71 , \P78:71 , \G78:71 );

  wire \P78:63 , \G78:63 ;

  PijGij \78:63 (\P78:71 , \P70:63 , \G78:71 , \G70:63 , \P78:63 , \G78:63 );

  wire \G78:-1 ;

  Gij \78:-1 (\P78:63 , \G78:63 , \G62:-1 , \G78:-1 );

  Sum s79(\G78:-1 , A[79], B[79], S[79]);

  wire \P79:63 , \G79:63 ;

  PijGij \79:63 (P[79], \P78:63 , G[79], \G78:63 , \P79:63 , \G79:63 );

  wire \G79:-1 ;

  Gij \79:-1 (\P79:63 , \G79:63 , \G62:-1 , \G79:-1 );

  Sum s80(\G79:-1 , A[80], B[80], S[80]);

  wire \P80:79 , \G80:79 ;

  PijGij \80:79 (P[80], P[79], G[80], G[79], \P80:79 , \G80:79 );

  wire \P80:63 , \G80:63 ;

  PijGij \80:63 (\P80:79 , \P78:63 , \G80:79 , \G78:63 , \P80:63 , \G80:63 );

  wire \G80:-1 ;

  Gij \80:-1 (\P80:63 , \G80:63 , \G62:-1 , \G80:-1 );

  Sum s81(\G80:-1 , A[81], B[81], S[81]);

  wire \P81:79 , \G81:79 ;

  PijGij \81:79 (P[81], \P80:79 , G[81], \G80:79 , \P81:79 , \G81:79 );

  wire \P81:63 , \G81:63 ;

  PijGij \81:63 (\P81:79 , \P78:63 , \G81:79 , \G78:63 , \P81:63 , \G81:63 );

  wire \G81:-1 ;

  Gij \81:-1 (\P81:63 , \G81:63 , \G62:-1 , \G81:-1 );

  Sum s82(\G81:-1 , A[82], B[82], S[82]);

  wire \P82:81 , \G82:81 ;

  PijGij \82:81 (P[82], P[81], G[82], G[81], \P82:81 , \G82:81 );

  wire \P82:79 , \G82:79 ;

  PijGij \82:79 (\P82:81 , \P80:79 , \G82:81 , \G80:79 , \P82:79 , \G82:79 );

  wire \P82:63 , \G82:63 ;

  PijGij \82:63 (\P82:79 , \P78:63 , \G82:79 , \G78:63 , \P82:63 , \G82:63 );

  wire \G82:-1 ;

  Gij \82:-1 (\P82:63 , \G82:63 , \G62:-1 , \G82:-1 );

  Sum s83(\G82:-1 , A[83], B[83], S[83]);

  wire \P83:79 , \G83:79 ;

  PijGij \83:79 (P[83], \P82:79 , G[83], \G82:79 , \P83:79 , \G83:79 );

  wire \P83:63 , \G83:63 ;

  PijGij \83:63 (\P83:79 , \P78:63 , \G83:79 , \G78:63 , \P83:63 , \G83:63 );

  wire \G83:-1 ;

  Gij \83:-1 (\P83:63 , \G83:63 , \G62:-1 , \G83:-1 );

  Sum s84(\G83:-1 , A[84], B[84], S[84]);

  wire \P84:83 , \G84:83 ;

  PijGij \84:83 (P[84], P[83], G[84], G[83], \P84:83 , \G84:83 );

  wire \P84:79 , \G84:79 ;

  PijGij \84:79 (\P84:83 , \P82:79 , \G84:83 , \G82:79 , \P84:79 , \G84:79 );

  wire \P84:63 , \G84:63 ;

  PijGij \84:63 (\P84:79 , \P78:63 , \G84:79 , \G78:63 , \P84:63 , \G84:63 );

  wire \G84:-1 ;

  Gij \84:-1 (\P84:63 , \G84:63 , \G62:-1 , \G84:-1 );

  Sum s85(\G84:-1 , A[85], B[85], S[85]);

  wire \P85:83 , \G85:83 ;

  PijGij \85:83 (P[85], \P84:83 , G[85], \G84:83 , \P85:83 , \G85:83 );

  wire \P85:79 , \G85:79 ;

  PijGij \85:79 (\P85:83 , \P82:79 , \G85:83 , \G82:79 , \P85:79 , \G85:79 );

  wire \P85:63 , \G85:63 ;

  PijGij \85:63 (\P85:79 , \P78:63 , \G85:79 , \G78:63 , \P85:63 , \G85:63 );

  wire \G85:-1 ;

  Gij \85:-1 (\P85:63 , \G85:63 , \G62:-1 , \G85:-1 );

  Sum s86(\G85:-1 , A[86], B[86], S[86]);

  wire \P86:85 , \G86:85 ;

  PijGij \86:85 (P[86], P[85], G[86], G[85], \P86:85 , \G86:85 );

  wire \P86:83 , \G86:83 ;

  PijGij \86:83 (\P86:85 , \P84:83 , \G86:85 , \G84:83 , \P86:83 , \G86:83 );

  wire \P86:79 , \G86:79 ;

  PijGij \86:79 (\P86:83 , \P82:79 , \G86:83 , \G82:79 , \P86:79 , \G86:79 );

  wire \P86:63 , \G86:63 ;

  PijGij \86:63 (\P86:79 , \P78:63 , \G86:79 , \G78:63 , \P86:63 , \G86:63 );

  wire \G86:-1 ;

  Gij \86:-1 (\P86:63 , \G86:63 , \G62:-1 , \G86:-1 );

  Sum s87(\G86:-1 , A[87], B[87], S[87]);

  wire \P87:79 , \G87:79 ;

  PijGij \87:79 (P[87], \P86:79 , G[87], \G86:79 , \P87:79 , \G87:79 );

  wire \P87:63 , \G87:63 ;

  PijGij \87:63 (\P87:79 , \P78:63 , \G87:79 , \G78:63 , \P87:63 , \G87:63 );

  wire \G87:-1 ;

  Gij \87:-1 (\P87:63 , \G87:63 , \G62:-1 , \G87:-1 );

  Sum s88(\G87:-1 , A[88], B[88], S[88]);

  wire \P88:87 , \G88:87 ;

  PijGij \88:87 (P[88], P[87], G[88], G[87], \P88:87 , \G88:87 );

  wire \P88:79 , \G88:79 ;

  PijGij \88:79 (\P88:87 , \P86:79 , \G88:87 , \G86:79 , \P88:79 , \G88:79 );

  wire \P88:63 , \G88:63 ;

  PijGij \88:63 (\P88:79 , \P78:63 , \G88:79 , \G78:63 , \P88:63 , \G88:63 );

  wire \G88:-1 ;

  Gij \88:-1 (\P88:63 , \G88:63 , \G62:-1 , \G88:-1 );

  Sum s89(\G88:-1 , A[89], B[89], S[89]);

  wire \P89:87 , \G89:87 ;

  PijGij \89:87 (P[89], \P88:87 , G[89], \G88:87 , \P89:87 , \G89:87 );

  wire \P89:79 , \G89:79 ;

  PijGij \89:79 (\P89:87 , \P86:79 , \G89:87 , \G86:79 , \P89:79 , \G89:79 );

  wire \P89:63 , \G89:63 ;

  PijGij \89:63 (\P89:79 , \P78:63 , \G89:79 , \G78:63 , \P89:63 , \G89:63 );

  wire \G89:-1 ;

  Gij \89:-1 (\P89:63 , \G89:63 , \G62:-1 , \G89:-1 );

  Sum s90(\G89:-1 , A[90], B[90], S[90]);

  wire \P90:89 , \G90:89 ;

  PijGij \90:89 (P[90], P[89], G[90], G[89], \P90:89 , \G90:89 );

  wire \P90:87 , \G90:87 ;

  PijGij \90:87 (\P90:89 , \P88:87 , \G90:89 , \G88:87 , \P90:87 , \G90:87 );

  wire \P90:79 , \G90:79 ;

  PijGij \90:79 (\P90:87 , \P86:79 , \G90:87 , \G86:79 , \P90:79 , \G90:79 );

  wire \P90:63 , \G90:63 ;

  PijGij \90:63 (\P90:79 , \P78:63 , \G90:79 , \G78:63 , \P90:63 , \G90:63 );

  wire \G90:-1 ;

  Gij \90:-1 (\P90:63 , \G90:63 , \G62:-1 , \G90:-1 );

  Sum s91(\G90:-1 , A[91], B[91], S[91]);

  wire \P91:87 , \G91:87 ;

  PijGij \91:87 (P[91], \P90:87 , G[91], \G90:87 , \P91:87 , \G91:87 );

  wire \P91:79 , \G91:79 ;

  PijGij \91:79 (\P91:87 , \P86:79 , \G91:87 , \G86:79 , \P91:79 , \G91:79 );

  wire \P91:63 , \G91:63 ;

  PijGij \91:63 (\P91:79 , \P78:63 , \G91:79 , \G78:63 , \P91:63 , \G91:63 );

  wire \G91:-1 ;

  Gij \91:-1 (\P91:63 , \G91:63 , \G62:-1 , \G91:-1 );

  Sum s92(\G91:-1 , A[92], B[92], S[92]);

  wire \P92:91 , \G92:91 ;

  PijGij \92:91 (P[92], P[91], G[92], G[91], \P92:91 , \G92:91 );

  wire \P92:87 , \G92:87 ;

  PijGij \92:87 (\P92:91 , \P90:87 , \G92:91 , \G90:87 , \P92:87 , \G92:87 );

  wire \P92:79 , \G92:79 ;

  PijGij \92:79 (\P92:87 , \P86:79 , \G92:87 , \G86:79 , \P92:79 , \G92:79 );

  wire \P92:63 , \G92:63 ;

  PijGij \92:63 (\P92:79 , \P78:63 , \G92:79 , \G78:63 , \P92:63 , \G92:63 );

  wire \G92:-1 ;

  Gij \92:-1 (\P92:63 , \G92:63 , \G62:-1 , \G92:-1 );

  Sum s93(\G92:-1 , A[93], B[93], S[93]);

  wire \P93:91 , \G93:91 ;

  PijGij \93:91 (P[93], \P92:91 , G[93], \G92:91 , \P93:91 , \G93:91 );

  wire \P93:87 , \G93:87 ;

  PijGij \93:87 (\P93:91 , \P90:87 , \G93:91 , \G90:87 , \P93:87 , \G93:87 );

  wire \P93:79 , \G93:79 ;

  PijGij \93:79 (\P93:87 , \P86:79 , \G93:87 , \G86:79 , \P93:79 , \G93:79 );

  wire \P93:63 , \G93:63 ;

  PijGij \93:63 (\P93:79 , \P78:63 , \G93:79 , \G78:63 , \P93:63 , \G93:63 );

  wire \G93:-1 ;

  Gij \93:-1 (\P93:63 , \G93:63 , \G62:-1 , \G93:-1 );

  Sum s94(\G93:-1 , A[94], B[94], S[94]);

  wire \P94:93 , \G94:93 ;

  PijGij \94:93 (P[94], P[93], G[94], G[93], \P94:93 , \G94:93 );

  wire \P94:91 , \G94:91 ;

  PijGij \94:91 (\P94:93 , \P92:91 , \G94:93 , \G92:91 , \P94:91 , \G94:91 );

  wire \P94:87 , \G94:87 ;

  PijGij \94:87 (\P94:91 , \P90:87 , \G94:91 , \G90:87 , \P94:87 , \G94:87 );

  wire \P94:79 , \G94:79 ;

  PijGij \94:79 (\P94:87 , \P86:79 , \G94:87 , \G86:79 , \P94:79 , \G94:79 );

  wire \P94:63 , \G94:63 ;

  PijGij \94:63 (\P94:79 , \P78:63 , \G94:79 , \G78:63 , \P94:63 , \G94:63 );

  wire \G94:-1 ;

  Gij \94:-1 (\P94:63 , \G94:63 , \G62:-1 , \G94:-1 );

  Sum s95(\G94:-1 , A[95], B[95], S[95]);

  wire \P95:63 , \G95:63 ;

  PijGij \95:63 (P[95], \P94:63 , G[95], \G94:63 , \P95:63 , \G95:63 );

  wire \G95:-1 ;

  Gij \95:-1 (\P95:63 , \G95:63 , \G62:-1 , \G95:-1 );

  Sum s96(\G95:-1 , A[96], B[96], S[96]);

  wire \P96:95 , \G96:95 ;

  PijGij \96:95 (P[96], P[95], G[96], G[95], \P96:95 , \G96:95 );

  wire \P96:63 , \G96:63 ;

  PijGij \96:63 (\P96:95 , \P94:63 , \G96:95 , \G94:63 , \P96:63 , \G96:63 );

  wire \G96:-1 ;

  Gij \96:-1 (\P96:63 , \G96:63 , \G62:-1 , \G96:-1 );

  Sum s97(\G96:-1 , A[97], B[97], S[97]);

  wire \P97:95 , \G97:95 ;

  PijGij \97:95 (P[97], \P96:95 , G[97], \G96:95 , \P97:95 , \G97:95 );

  wire \P97:63 , \G97:63 ;

  PijGij \97:63 (\P97:95 , \P94:63 , \G97:95 , \G94:63 , \P97:63 , \G97:63 );

  wire \G97:-1 ;

  Gij \97:-1 (\P97:63 , \G97:63 , \G62:-1 , \G97:-1 );

  Sum s98(\G97:-1 , A[98], B[98], S[98]);

  wire \P98:97 , \G98:97 ;

  PijGij \98:97 (P[98], P[97], G[98], G[97], \P98:97 , \G98:97 );

  wire \P98:95 , \G98:95 ;

  PijGij \98:95 (\P98:97 , \P96:95 , \G98:97 , \G96:95 , \P98:95 , \G98:95 );

  wire \P98:63 , \G98:63 ;

  PijGij \98:63 (\P98:95 , \P94:63 , \G98:95 , \G94:63 , \P98:63 , \G98:63 );

  wire \G98:-1 ;

  Gij \98:-1 (\P98:63 , \G98:63 , \G62:-1 , \G98:-1 );

  Sum s99(\G98:-1 , A[99], B[99], S[99]);

  wire \P99:95 , \G99:95 ;

  PijGij \99:95 (P[99], \P98:95 , G[99], \G98:95 , \P99:95 , \G99:95 );

  wire \P99:63 , \G99:63 ;

  PijGij \99:63 (\P99:95 , \P94:63 , \G99:95 , \G94:63 , \P99:63 , \G99:63 );

  wire \G99:-1 ;

  Gij \99:-1 (\P99:63 , \G99:63 , \G62:-1 , \G99:-1 );

  Sum s100(\G99:-1 , A[100], B[100], S[100]);

  wire \P100:99 , \G100:99 ;

  PijGij \100:99 (P[100], P[99], G[100], G[99], \P100:99 , \G100:99 );

  wire \P100:95 , \G100:95 ;

  PijGij \100:95 (\P100:99 , \P98:95 , \G100:99 , \G98:95 , \P100:95 , \G100:95 );

  wire \P100:63 , \G100:63 ;

  PijGij \100:63 (\P100:95 , \P94:63 , \G100:95 , \G94:63 , \P100:63 , \G100:63 );

  wire \G100:-1 ;

  Gij \100:-1 (\P100:63 , \G100:63 , \G62:-1 , \G100:-1 );

  Sum s101(\G100:-1 , A[101], B[101], S[101]);

  wire \P101:99 , \G101:99 ;

  PijGij \101:99 (P[101], \P100:99 , G[101], \G100:99 , \P101:99 , \G101:99 );

  wire \P101:95 , \G101:95 ;

  PijGij \101:95 (\P101:99 , \P98:95 , \G101:99 , \G98:95 , \P101:95 , \G101:95 );

  wire \P101:63 , \G101:63 ;

  PijGij \101:63 (\P101:95 , \P94:63 , \G101:95 , \G94:63 , \P101:63 , \G101:63 );

  wire \G101:-1 ;

  Gij \101:-1 (\P101:63 , \G101:63 , \G62:-1 , \G101:-1 );

  Sum s102(\G101:-1 , A[102], B[102], S[102]);

  wire \P102:101 , \G102:101 ;

  PijGij \102:101 (P[102], P[101], G[102], G[101], \P102:101 , \G102:101 );

  wire \P102:99 , \G102:99 ;

  PijGij \102:99 (\P102:101 , \P100:99 , \G102:101 , \G100:99 , \P102:99 , \G102:99 );

  wire \P102:95 , \G102:95 ;

  PijGij \102:95 (\P102:99 , \P98:95 , \G102:99 , \G98:95 , \P102:95 , \G102:95 );

  wire \P102:63 , \G102:63 ;

  PijGij \102:63 (\P102:95 , \P94:63 , \G102:95 , \G94:63 , \P102:63 , \G102:63 );

  wire \G102:-1 ;

  Gij \102:-1 (\P102:63 , \G102:63 , \G62:-1 , \G102:-1 );

  Sum s103(\G102:-1 , A[103], B[103], S[103]);

  wire \P103:95 , \G103:95 ;

  PijGij \103:95 (P[103], \P102:95 , G[103], \G102:95 , \P103:95 , \G103:95 );

  wire \P103:63 , \G103:63 ;

  PijGij \103:63 (\P103:95 , \P94:63 , \G103:95 , \G94:63 , \P103:63 , \G103:63 );

  wire \G103:-1 ;

  Gij \103:-1 (\P103:63 , \G103:63 , \G62:-1 , \G103:-1 );

  Sum s104(\G103:-1 , A[104], B[104], S[104]);

  wire \P104:103 , \G104:103 ;

  PijGij \104:103 (P[104], P[103], G[104], G[103], \P104:103 , \G104:103 );

  wire \P104:95 , \G104:95 ;

  PijGij \104:95 (\P104:103 , \P102:95 , \G104:103 , \G102:95 , \P104:95 , \G104:95 );

  wire \P104:63 , \G104:63 ;

  PijGij \104:63 (\P104:95 , \P94:63 , \G104:95 , \G94:63 , \P104:63 , \G104:63 );

  wire \G104:-1 ;

  Gij \104:-1 (\P104:63 , \G104:63 , \G62:-1 , \G104:-1 );

  Sum s105(\G104:-1 , A[105], B[105], S[105]);

  wire \P105:103 , \G105:103 ;

  PijGij \105:103 (P[105], \P104:103 , G[105], \G104:103 , \P105:103 , \G105:103 );

  wire \P105:95 , \G105:95 ;

  PijGij \105:95 (\P105:103 , \P102:95 , \G105:103 , \G102:95 , \P105:95 , \G105:95 );

  wire \P105:63 , \G105:63 ;

  PijGij \105:63 (\P105:95 , \P94:63 , \G105:95 , \G94:63 , \P105:63 , \G105:63 );

  wire \G105:-1 ;

  Gij \105:-1 (\P105:63 , \G105:63 , \G62:-1 , \G105:-1 );

  Sum s106(\G105:-1 , A[106], B[106], S[106]);

  wire \P106:105 , \G106:105 ;

  PijGij \106:105 (P[106], P[105], G[106], G[105], \P106:105 , \G106:105 );

  wire \P106:103 , \G106:103 ;

  PijGij \106:103 (\P106:105 , \P104:103 , \G106:105 , \G104:103 , \P106:103 , \G106:103 );

  wire \P106:95 , \G106:95 ;

  PijGij \106:95 (\P106:103 , \P102:95 , \G106:103 , \G102:95 , \P106:95 , \G106:95 );

  wire \P106:63 , \G106:63 ;

  PijGij \106:63 (\P106:95 , \P94:63 , \G106:95 , \G94:63 , \P106:63 , \G106:63 );

  wire \G106:-1 ;

  Gij \106:-1 (\P106:63 , \G106:63 , \G62:-1 , \G106:-1 );

  Sum s107(\G106:-1 , A[107], B[107], S[107]);

  wire \P107:103 , \G107:103 ;

  PijGij \107:103 (P[107], \P106:103 , G[107], \G106:103 , \P107:103 , \G107:103 );

  wire \P107:95 , \G107:95 ;

  PijGij \107:95 (\P107:103 , \P102:95 , \G107:103 , \G102:95 , \P107:95 , \G107:95 );

  wire \P107:63 , \G107:63 ;

  PijGij \107:63 (\P107:95 , \P94:63 , \G107:95 , \G94:63 , \P107:63 , \G107:63 );

  wire \G107:-1 ;

  Gij \107:-1 (\P107:63 , \G107:63 , \G62:-1 , \G107:-1 );

  Sum s108(\G107:-1 , A[108], B[108], S[108]);

  wire \P108:107 , \G108:107 ;

  PijGij \108:107 (P[108], P[107], G[108], G[107], \P108:107 , \G108:107 );

  wire \P108:103 , \G108:103 ;

  PijGij \108:103 (\P108:107 , \P106:103 , \G108:107 , \G106:103 , \P108:103 , \G108:103 );

  wire \P108:95 , \G108:95 ;

  PijGij \108:95 (\P108:103 , \P102:95 , \G108:103 , \G102:95 , \P108:95 , \G108:95 );

  wire \P108:63 , \G108:63 ;

  PijGij \108:63 (\P108:95 , \P94:63 , \G108:95 , \G94:63 , \P108:63 , \G108:63 );

  wire \G108:-1 ;

  Gij \108:-1 (\P108:63 , \G108:63 , \G62:-1 , \G108:-1 );

  Sum s109(\G108:-1 , A[109], B[109], S[109]);

  wire \P109:107 , \G109:107 ;

  PijGij \109:107 (P[109], \P108:107 , G[109], \G108:107 , \P109:107 , \G109:107 );

  wire \P109:103 , \G109:103 ;

  PijGij \109:103 (\P109:107 , \P106:103 , \G109:107 , \G106:103 , \P109:103 , \G109:103 );

  wire \P109:95 , \G109:95 ;

  PijGij \109:95 (\P109:103 , \P102:95 , \G109:103 , \G102:95 , \P109:95 , \G109:95 );

  wire \P109:63 , \G109:63 ;

  PijGij \109:63 (\P109:95 , \P94:63 , \G109:95 , \G94:63 , \P109:63 , \G109:63 );

  wire \G109:-1 ;

  Gij \109:-1 (\P109:63 , \G109:63 , \G62:-1 , \G109:-1 );

  Sum s110(\G109:-1 , A[110], B[110], S[110]);

  wire \P110:109 , \G110:109 ;

  PijGij \110:109 (P[110], P[109], G[110], G[109], \P110:109 , \G110:109 );

  wire \P110:107 , \G110:107 ;

  PijGij \110:107 (\P110:109 , \P108:107 , \G110:109 , \G108:107 , \P110:107 , \G110:107 );

  wire \P110:103 , \G110:103 ;

  PijGij \110:103 (\P110:107 , \P106:103 , \G110:107 , \G106:103 , \P110:103 , \G110:103 );

  wire \P110:95 , \G110:95 ;

  PijGij \110:95 (\P110:103 , \P102:95 , \G110:103 , \G102:95 , \P110:95 , \G110:95 );

  wire \P110:63 , \G110:63 ;

  PijGij \110:63 (\P110:95 , \P94:63 , \G110:95 , \G94:63 , \P110:63 , \G110:63 );

  wire \G110:-1 ;

  Gij \110:-1 (\P110:63 , \G110:63 , \G62:-1 , \G110:-1 );

  Sum s111(\G110:-1 , A[111], B[111], S[111]);

  wire \P111:95 , \G111:95 ;

  PijGij \111:95 (P[111], \P110:95 , G[111], \G110:95 , \P111:95 , \G111:95 );

  wire \P111:63 , \G111:63 ;

  PijGij \111:63 (\P111:95 , \P94:63 , \G111:95 , \G94:63 , \P111:63 , \G111:63 );

  wire \G111:-1 ;

  Gij \111:-1 (\P111:63 , \G111:63 , \G62:-1 , \G111:-1 );

  Sum s112(\G111:-1 , A[112], B[112], S[112]);

  wire \P112:111 , \G112:111 ;

  PijGij \112:111 (P[112], P[111], G[112], G[111], \P112:111 , \G112:111 );

  wire \P112:95 , \G112:95 ;

  PijGij \112:95 (\P112:111 , \P110:95 , \G112:111 , \G110:95 , \P112:95 , \G112:95 );

  wire \P112:63 , \G112:63 ;

  PijGij \112:63 (\P112:95 , \P94:63 , \G112:95 , \G94:63 , \P112:63 , \G112:63 );

  wire \G112:-1 ;

  Gij \112:-1 (\P112:63 , \G112:63 , \G62:-1 , \G112:-1 );

  Sum s113(\G112:-1 , A[113], B[113], S[113]);

  wire \P113:111 , \G113:111 ;

  PijGij \113:111 (P[113], \P112:111 , G[113], \G112:111 , \P113:111 , \G113:111 );

  wire \P113:95 , \G113:95 ;

  PijGij \113:95 (\P113:111 , \P110:95 , \G113:111 , \G110:95 , \P113:95 , \G113:95 );

  wire \P113:63 , \G113:63 ;

  PijGij \113:63 (\P113:95 , \P94:63 , \G113:95 , \G94:63 , \P113:63 , \G113:63 );

  wire \G113:-1 ;

  Gij \113:-1 (\P113:63 , \G113:63 , \G62:-1 , \G113:-1 );

  Sum s114(\G113:-1 , A[114], B[114], S[114]);

  wire \P114:113 , \G114:113 ;

  PijGij \114:113 (P[114], P[113], G[114], G[113], \P114:113 , \G114:113 );

  wire \P114:111 , \G114:111 ;

  PijGij \114:111 (\P114:113 , \P112:111 , \G114:113 , \G112:111 , \P114:111 , \G114:111 );

  wire \P114:95 , \G114:95 ;

  PijGij \114:95 (\P114:111 , \P110:95 , \G114:111 , \G110:95 , \P114:95 , \G114:95 );

  wire \P114:63 , \G114:63 ;

  PijGij \114:63 (\P114:95 , \P94:63 , \G114:95 , \G94:63 , \P114:63 , \G114:63 );

  wire \G114:-1 ;

  Gij \114:-1 (\P114:63 , \G114:63 , \G62:-1 , \G114:-1 );

  Sum s115(\G114:-1 , A[115], B[115], S[115]);

  wire \P115:111 , \G115:111 ;

  PijGij \115:111 (P[115], \P114:111 , G[115], \G114:111 , \P115:111 , \G115:111 );

  wire \P115:95 , \G115:95 ;

  PijGij \115:95 (\P115:111 , \P110:95 , \G115:111 , \G110:95 , \P115:95 , \G115:95 );

  wire \P115:63 , \G115:63 ;

  PijGij \115:63 (\P115:95 , \P94:63 , \G115:95 , \G94:63 , \P115:63 , \G115:63 );

  wire \G115:-1 ;

  Gij \115:-1 (\P115:63 , \G115:63 , \G62:-1 , \G115:-1 );

  Sum s116(\G115:-1 , A[116], B[116], S[116]);

  wire \P116:115 , \G116:115 ;

  PijGij \116:115 (P[116], P[115], G[116], G[115], \P116:115 , \G116:115 );

  wire \P116:111 , \G116:111 ;

  PijGij \116:111 (\P116:115 , \P114:111 , \G116:115 , \G114:111 , \P116:111 , \G116:111 );

  wire \P116:95 , \G116:95 ;

  PijGij \116:95 (\P116:111 , \P110:95 , \G116:111 , \G110:95 , \P116:95 , \G116:95 );

  wire \P116:63 , \G116:63 ;

  PijGij \116:63 (\P116:95 , \P94:63 , \G116:95 , \G94:63 , \P116:63 , \G116:63 );

  wire \G116:-1 ;

  Gij \116:-1 (\P116:63 , \G116:63 , \G62:-1 , \G116:-1 );

  Sum s117(\G116:-1 , A[117], B[117], S[117]);

  wire \P117:115 , \G117:115 ;

  PijGij \117:115 (P[117], \P116:115 , G[117], \G116:115 , \P117:115 , \G117:115 );

  wire \P117:111 , \G117:111 ;

  PijGij \117:111 (\P117:115 , \P114:111 , \G117:115 , \G114:111 , \P117:111 , \G117:111 );

  wire \P117:95 , \G117:95 ;

  PijGij \117:95 (\P117:111 , \P110:95 , \G117:111 , \G110:95 , \P117:95 , \G117:95 );

  wire \P117:63 , \G117:63 ;

  PijGij \117:63 (\P117:95 , \P94:63 , \G117:95 , \G94:63 , \P117:63 , \G117:63 );

  wire \G117:-1 ;

  Gij \117:-1 (\P117:63 , \G117:63 , \G62:-1 , \G117:-1 );

  Sum s118(\G117:-1 , A[118], B[118], S[118]);

  wire \P118:117 , \G118:117 ;

  PijGij \118:117 (P[118], P[117], G[118], G[117], \P118:117 , \G118:117 );

  wire \P118:115 , \G118:115 ;

  PijGij \118:115 (\P118:117 , \P116:115 , \G118:117 , \G116:115 , \P118:115 , \G118:115 );

  wire \P118:111 , \G118:111 ;

  PijGij \118:111 (\P118:115 , \P114:111 , \G118:115 , \G114:111 , \P118:111 , \G118:111 );

  wire \P118:95 , \G118:95 ;

  PijGij \118:95 (\P118:111 , \P110:95 , \G118:111 , \G110:95 , \P118:95 , \G118:95 );

  wire \P118:63 , \G118:63 ;

  PijGij \118:63 (\P118:95 , \P94:63 , \G118:95 , \G94:63 , \P118:63 , \G118:63 );

  wire \G118:-1 ;

  Gij \118:-1 (\P118:63 , \G118:63 , \G62:-1 , \G118:-1 );

  Sum s119(\G118:-1 , A[119], B[119], S[119]);

  wire \P119:111 , \G119:111 ;

  PijGij \119:111 (P[119], \P118:111 , G[119], \G118:111 , \P119:111 , \G119:111 );

  wire \P119:95 , \G119:95 ;

  PijGij \119:95 (\P119:111 , \P110:95 , \G119:111 , \G110:95 , \P119:95 , \G119:95 );

  wire \P119:63 , \G119:63 ;

  PijGij \119:63 (\P119:95 , \P94:63 , \G119:95 , \G94:63 , \P119:63 , \G119:63 );

  wire \G119:-1 ;

  Gij \119:-1 (\P119:63 , \G119:63 , \G62:-1 , \G119:-1 );

  Sum s120(\G119:-1 , A[120], B[120], S[120]);

  wire \P120:119 , \G120:119 ;

  PijGij \120:119 (P[120], P[119], G[120], G[119], \P120:119 , \G120:119 );

  wire \P120:111 , \G120:111 ;

  PijGij \120:111 (\P120:119 , \P118:111 , \G120:119 , \G118:111 , \P120:111 , \G120:111 );

  wire \P120:95 , \G120:95 ;

  PijGij \120:95 (\P120:111 , \P110:95 , \G120:111 , \G110:95 , \P120:95 , \G120:95 );

  wire \P120:63 , \G120:63 ;

  PijGij \120:63 (\P120:95 , \P94:63 , \G120:95 , \G94:63 , \P120:63 , \G120:63 );

  wire \G120:-1 ;

  Gij \120:-1 (\P120:63 , \G120:63 , \G62:-1 , \G120:-1 );

  Sum s121(\G120:-1 , A[121], B[121], S[121]);

  wire \P121:119 , \G121:119 ;

  PijGij \121:119 (P[121], \P120:119 , G[121], \G120:119 , \P121:119 , \G121:119 );

  wire \P121:111 , \G121:111 ;

  PijGij \121:111 (\P121:119 , \P118:111 , \G121:119 , \G118:111 , \P121:111 , \G121:111 );

  wire \P121:95 , \G121:95 ;

  PijGij \121:95 (\P121:111 , \P110:95 , \G121:111 , \G110:95 , \P121:95 , \G121:95 );

  wire \P121:63 , \G121:63 ;

  PijGij \121:63 (\P121:95 , \P94:63 , \G121:95 , \G94:63 , \P121:63 , \G121:63 );

  wire \G121:-1 ;

  Gij \121:-1 (\P121:63 , \G121:63 , \G62:-1 , \G121:-1 );

  Sum s122(\G121:-1 , A[122], B[122], S[122]);

  wire \P122:121 , \G122:121 ;

  PijGij \122:121 (P[122], P[121], G[122], G[121], \P122:121 , \G122:121 );

  wire \P122:119 , \G122:119 ;

  PijGij \122:119 (\P122:121 , \P120:119 , \G122:121 , \G120:119 , \P122:119 , \G122:119 );

  wire \P122:111 , \G122:111 ;

  PijGij \122:111 (\P122:119 , \P118:111 , \G122:119 , \G118:111 , \P122:111 , \G122:111 );

  wire \P122:95 , \G122:95 ;

  PijGij \122:95 (\P122:111 , \P110:95 , \G122:111 , \G110:95 , \P122:95 , \G122:95 );

  wire \P122:63 , \G122:63 ;

  PijGij \122:63 (\P122:95 , \P94:63 , \G122:95 , \G94:63 , \P122:63 , \G122:63 );

  wire \G122:-1 ;

  Gij \122:-1 (\P122:63 , \G122:63 , \G62:-1 , \G122:-1 );

  Sum s123(\G122:-1 , A[123], B[123], S[123]);

  wire \P123:119 , \G123:119 ;

  PijGij \123:119 (P[123], \P122:119 , G[123], \G122:119 , \P123:119 , \G123:119 );

  wire \P123:111 , \G123:111 ;

  PijGij \123:111 (\P123:119 , \P118:111 , \G123:119 , \G118:111 , \P123:111 , \G123:111 );

  wire \P123:95 , \G123:95 ;

  PijGij \123:95 (\P123:111 , \P110:95 , \G123:111 , \G110:95 , \P123:95 , \G123:95 );

  wire \P123:63 , \G123:63 ;

  PijGij \123:63 (\P123:95 , \P94:63 , \G123:95 , \G94:63 , \P123:63 , \G123:63 );

  wire \G123:-1 ;

  Gij \123:-1 (\P123:63 , \G123:63 , \G62:-1 , \G123:-1 );

  Sum s124(\G123:-1 , A[124], B[124], S[124]);

  wire \P124:123 , \G124:123 ;

  PijGij \124:123 (P[124], P[123], G[124], G[123], \P124:123 , \G124:123 );

  wire \P124:119 , \G124:119 ;

  PijGij \124:119 (\P124:123 , \P122:119 , \G124:123 , \G122:119 , \P124:119 , \G124:119 );

  wire \P124:111 , \G124:111 ;

  PijGij \124:111 (\P124:119 , \P118:111 , \G124:119 , \G118:111 , \P124:111 , \G124:111 );

  wire \P124:95 , \G124:95 ;

  PijGij \124:95 (\P124:111 , \P110:95 , \G124:111 , \G110:95 , \P124:95 , \G124:95 );

  wire \P124:63 , \G124:63 ;

  PijGij \124:63 (\P124:95 , \P94:63 , \G124:95 , \G94:63 , \P124:63 , \G124:63 );

  wire \G124:-1 ;

  Gij \124:-1 (\P124:63 , \G124:63 , \G62:-1 , \G124:-1 );

  Sum s125(\G124:-1 , A[125], B[125], S[125]);

  wire \P125:123 , \G125:123 ;

  PijGij \125:123 (P[125], \P124:123 , G[125], \G124:123 , \P125:123 , \G125:123 );

  wire \P125:119 , \G125:119 ;

  PijGij \125:119 (\P125:123 , \P122:119 , \G125:123 , \G122:119 , \P125:119 , \G125:119 );

  wire \P125:111 , \G125:111 ;

  PijGij \125:111 (\P125:119 , \P118:111 , \G125:119 , \G118:111 , \P125:111 , \G125:111 );

  wire \P125:95 , \G125:95 ;

  PijGij \125:95 (\P125:111 , \P110:95 , \G125:111 , \G110:95 , \P125:95 , \G125:95 );

  wire \P125:63 , \G125:63 ;

  PijGij \125:63 (\P125:95 , \P94:63 , \G125:95 , \G94:63 , \P125:63 , \G125:63 );

  wire \G125:-1 ;

  Gij \125:-1 (\P125:63 , \G125:63 , \G62:-1 , \G125:-1 );

  Sum s126(\G125:-1 , A[126], B[126], S[126]);

  wire \P126:125 , \G126:125 ;

  PijGij \126:125 (P[126], P[125], G[126], G[125], \P126:125 , \G126:125 );

  wire \P126:123 , \G126:123 ;

  PijGij \126:123 (\P126:125 , \P124:123 , \G126:125 , \G124:123 , \P126:123 , \G126:123 );

  wire \P126:119 , \G126:119 ;

  PijGij \126:119 (\P126:123 , \P122:119 , \G126:123 , \G122:119 , \P126:119 , \G126:119 );

  wire \P126:111 , \G126:111 ;

  PijGij \126:111 (\P126:119 , \P118:111 , \G126:119 , \G118:111 , \P126:111 , \G126:111 );

  wire \P126:95 , \G126:95 ;

  PijGij \126:95 (\P126:111 , \P110:95 , \G126:111 , \G110:95 , \P126:95 , \G126:95 );

  wire \P126:63 , \G126:63 ;

  PijGij \126:63 (\P126:95 , \P94:63 , \G126:95 , \G94:63 , \P126:63 , \G126:63 );

  wire \G126:-1 ;

  Gij \126:-1 (\P126:63 , \G126:63 , \G62:-1 , \G126:-1 );

  Sum s127(\G126:-1 , A[127], B[127], S[127]);

  wire \G127:-1 ;

  Gij \127:-1 (P[127], G[127], \G126:-1 , \G127:-1 );

  Sum s128(\G127:-1 , A[128], B[128], S[128]);

  wire \P128:127 , \G128:127 ;

  PijGij \128:127 (P[128], P[127], G[128], G[127], \P128:127 , \G128:127 );

  wire \G128:-1 ;

  Gij \128:-1 (\P128:127 , \G128:127 , \G126:-1 , \G128:-1 );

  Sum s129(\G128:-1 , A[129], B[129], S[129]);

  wire \P129:127 , \G129:127 ;

  PijGij \129:127 (P[129], \P128:127 , G[129], \G128:127 , \P129:127 , \G129:127 );

  wire \G129:-1 ;

  Gij \129:-1 (\P129:127 , \G129:127 , \G126:-1 , \G129:-1 );

  Sum s130(\G129:-1 , A[130], B[130], S[130]);

  wire \P130:129 , \G130:129 ;

  PijGij \130:129 (P[130], P[129], G[130], G[129], \P130:129 , \G130:129 );

  wire \P130:127 , \G130:127 ;

  PijGij \130:127 (\P130:129 , \P128:127 , \G130:129 , \G128:127 , \P130:127 , \G130:127 );

  wire \G130:-1 ;

  Gij \130:-1 (\P130:127 , \G130:127 , \G126:-1 , \G130:-1 );

  Sum s131(\G130:-1 , A[131], B[131], S[131]);

  wire \P131:127 , \G131:127 ;

  PijGij \131:127 (P[131], \P130:127 , G[131], \G130:127 , \P131:127 , \G131:127 );

  wire \G131:-1 ;

  Gij \131:-1 (\P131:127 , \G131:127 , \G126:-1 , \G131:-1 );

  Sum s132(\G131:-1 , A[132], B[132], S[132]);

  wire \P132:131 , \G132:131 ;

  PijGij \132:131 (P[132], P[131], G[132], G[131], \P132:131 , \G132:131 );

  wire \P132:127 , \G132:127 ;

  PijGij \132:127 (\P132:131 , \P130:127 , \G132:131 , \G130:127 , \P132:127 , \G132:127 );

  wire \G132:-1 ;

  Gij \132:-1 (\P132:127 , \G132:127 , \G126:-1 , \G132:-1 );

  Sum s133(\G132:-1 , A[133], B[133], S[133]);

  wire \P133:131 , \G133:131 ;

  PijGij \133:131 (P[133], \P132:131 , G[133], \G132:131 , \P133:131 , \G133:131 );

  wire \P133:127 , \G133:127 ;

  PijGij \133:127 (\P133:131 , \P130:127 , \G133:131 , \G130:127 , \P133:127 , \G133:127 );

  wire \G133:-1 ;

  Gij \133:-1 (\P133:127 , \G133:127 , \G126:-1 , \G133:-1 );

  Sum s134(\G133:-1 , A[134], B[134], S[134]);

  wire \P134:133 , \G134:133 ;

  PijGij \134:133 (P[134], P[133], G[134], G[133], \P134:133 , \G134:133 );

  wire \P134:131 , \G134:131 ;

  PijGij \134:131 (\P134:133 , \P132:131 , \G134:133 , \G132:131 , \P134:131 , \G134:131 );

  wire \P134:127 , \G134:127 ;

  PijGij \134:127 (\P134:131 , \P130:127 , \G134:131 , \G130:127 , \P134:127 , \G134:127 );

  wire \G134:-1 ;

  Gij \134:-1 (\P134:127 , \G134:127 , \G126:-1 , \G134:-1 );

  Sum s135(\G134:-1 , A[135], B[135], S[135]);

  wire \P135:127 , \G135:127 ;

  PijGij \135:127 (P[135], \P134:127 , G[135], \G134:127 , \P135:127 , \G135:127 );

  wire \G135:-1 ;

  Gij \135:-1 (\P135:127 , \G135:127 , \G126:-1 , \G135:-1 );

  Sum s136(\G135:-1 , A[136], B[136], S[136]);

  wire \P136:135 , \G136:135 ;

  PijGij \136:135 (P[136], P[135], G[136], G[135], \P136:135 , \G136:135 );

  wire \P136:127 , \G136:127 ;

  PijGij \136:127 (\P136:135 , \P134:127 , \G136:135 , \G134:127 , \P136:127 , \G136:127 );

  wire \G136:-1 ;

  Gij \136:-1 (\P136:127 , \G136:127 , \G126:-1 , \G136:-1 );

  Sum s137(\G136:-1 , A[137], B[137], S[137]);

  wire \P137:135 , \G137:135 ;

  PijGij \137:135 (P[137], \P136:135 , G[137], \G136:135 , \P137:135 , \G137:135 );

  wire \P137:127 , \G137:127 ;

  PijGij \137:127 (\P137:135 , \P134:127 , \G137:135 , \G134:127 , \P137:127 , \G137:127 );

  wire \G137:-1 ;

  Gij \137:-1 (\P137:127 , \G137:127 , \G126:-1 , \G137:-1 );

  Sum s138(\G137:-1 , A[138], B[138], S[138]);

  wire \P138:137 , \G138:137 ;

  PijGij \138:137 (P[138], P[137], G[138], G[137], \P138:137 , \G138:137 );

  wire \P138:135 , \G138:135 ;

  PijGij \138:135 (\P138:137 , \P136:135 , \G138:137 , \G136:135 , \P138:135 , \G138:135 );

  wire \P138:127 , \G138:127 ;

  PijGij \138:127 (\P138:135 , \P134:127 , \G138:135 , \G134:127 , \P138:127 , \G138:127 );

  wire \G138:-1 ;

  Gij \138:-1 (\P138:127 , \G138:127 , \G126:-1 , \G138:-1 );

  Sum s139(\G138:-1 , A[139], B[139], S[139]);

  wire \P139:135 , \G139:135 ;

  PijGij \139:135 (P[139], \P138:135 , G[139], \G138:135 , \P139:135 , \G139:135 );

  wire \P139:127 , \G139:127 ;

  PijGij \139:127 (\P139:135 , \P134:127 , \G139:135 , \G134:127 , \P139:127 , \G139:127 );

  wire \G139:-1 ;

  Gij \139:-1 (\P139:127 , \G139:127 , \G126:-1 , \G139:-1 );

  Sum s140(\G139:-1 , A[140], B[140], S[140]);

  wire \P140:139 , \G140:139 ;

  PijGij \140:139 (P[140], P[139], G[140], G[139], \P140:139 , \G140:139 );

  wire \P140:135 , \G140:135 ;

  PijGij \140:135 (\P140:139 , \P138:135 , \G140:139 , \G138:135 , \P140:135 , \G140:135 );

  wire \P140:127 , \G140:127 ;

  PijGij \140:127 (\P140:135 , \P134:127 , \G140:135 , \G134:127 , \P140:127 , \G140:127 );

  wire \G140:-1 ;

  Gij \140:-1 (\P140:127 , \G140:127 , \G126:-1 , \G140:-1 );

  Sum s141(\G140:-1 , A[141], B[141], S[141]);

  wire \P141:139 , \G141:139 ;

  PijGij \141:139 (P[141], \P140:139 , G[141], \G140:139 , \P141:139 , \G141:139 );

  wire \P141:135 , \G141:135 ;

  PijGij \141:135 (\P141:139 , \P138:135 , \G141:139 , \G138:135 , \P141:135 , \G141:135 );

  wire \P141:127 , \G141:127 ;

  PijGij \141:127 (\P141:135 , \P134:127 , \G141:135 , \G134:127 , \P141:127 , \G141:127 );

  wire \G141:-1 ;

  Gij \141:-1 (\P141:127 , \G141:127 , \G126:-1 , \G141:-1 );

  Sum s142(\G141:-1 , A[142], B[142], S[142]);

  wire \P142:141 , \G142:141 ;

  PijGij \142:141 (P[142], P[141], G[142], G[141], \P142:141 , \G142:141 );

  wire \P142:139 , \G142:139 ;

  PijGij \142:139 (\P142:141 , \P140:139 , \G142:141 , \G140:139 , \P142:139 , \G142:139 );

  wire \P142:135 , \G142:135 ;

  PijGij \142:135 (\P142:139 , \P138:135 , \G142:139 , \G138:135 , \P142:135 , \G142:135 );

  wire \P142:127 , \G142:127 ;

  PijGij \142:127 (\P142:135 , \P134:127 , \G142:135 , \G134:127 , \P142:127 , \G142:127 );

  wire \G142:-1 ;

  Gij \142:-1 (\P142:127 , \G142:127 , \G126:-1 , \G142:-1 );

  Sum s143(\G142:-1 , A[143], B[143], S[143]);

  wire \P143:127 , \G143:127 ;

  PijGij \143:127 (P[143], \P142:127 , G[143], \G142:127 , \P143:127 , \G143:127 );

  wire \G143:-1 ;

  Gij \143:-1 (\P143:127 , \G143:127 , \G126:-1 , \G143:-1 );

  Sum s144(\G143:-1 , A[144], B[144], S[144]);

  wire \P144:143 , \G144:143 ;

  PijGij \144:143 (P[144], P[143], G[144], G[143], \P144:143 , \G144:143 );

  wire \P144:127 , \G144:127 ;

  PijGij \144:127 (\P144:143 , \P142:127 , \G144:143 , \G142:127 , \P144:127 , \G144:127 );

  wire \G144:-1 ;

  Gij \144:-1 (\P144:127 , \G144:127 , \G126:-1 , \G144:-1 );

  Sum s145(\G144:-1 , A[145], B[145], S[145]);

  wire \P145:143 , \G145:143 ;

  PijGij \145:143 (P[145], \P144:143 , G[145], \G144:143 , \P145:143 , \G145:143 );

  wire \P145:127 , \G145:127 ;

  PijGij \145:127 (\P145:143 , \P142:127 , \G145:143 , \G142:127 , \P145:127 , \G145:127 );

  wire \G145:-1 ;

  Gij \145:-1 (\P145:127 , \G145:127 , \G126:-1 , \G145:-1 );

  Sum s146(\G145:-1 , A[146], B[146], S[146]);

  wire \P146:145 , \G146:145 ;

  PijGij \146:145 (P[146], P[145], G[146], G[145], \P146:145 , \G146:145 );

  wire \P146:143 , \G146:143 ;

  PijGij \146:143 (\P146:145 , \P144:143 , \G146:145 , \G144:143 , \P146:143 , \G146:143 );

  wire \P146:127 , \G146:127 ;

  PijGij \146:127 (\P146:143 , \P142:127 , \G146:143 , \G142:127 , \P146:127 , \G146:127 );

  wire \G146:-1 ;

  Gij \146:-1 (\P146:127 , \G146:127 , \G126:-1 , \G146:-1 );

  Sum s147(\G146:-1 , A[147], B[147], S[147]);

  wire \P147:143 , \G147:143 ;

  PijGij \147:143 (P[147], \P146:143 , G[147], \G146:143 , \P147:143 , \G147:143 );

  wire \P147:127 , \G147:127 ;

  PijGij \147:127 (\P147:143 , \P142:127 , \G147:143 , \G142:127 , \P147:127 , \G147:127 );

  wire \G147:-1 ;

  Gij \147:-1 (\P147:127 , \G147:127 , \G126:-1 , \G147:-1 );

  Sum s148(\G147:-1 , A[148], B[148], S[148]);

  wire \P148:147 , \G148:147 ;

  PijGij \148:147 (P[148], P[147], G[148], G[147], \P148:147 , \G148:147 );

  wire \P148:143 , \G148:143 ;

  PijGij \148:143 (\P148:147 , \P146:143 , \G148:147 , \G146:143 , \P148:143 , \G148:143 );

  wire \P148:127 , \G148:127 ;

  PijGij \148:127 (\P148:143 , \P142:127 , \G148:143 , \G142:127 , \P148:127 , \G148:127 );

  wire \G148:-1 ;

  Gij \148:-1 (\P148:127 , \G148:127 , \G126:-1 , \G148:-1 );

  Sum s149(\G148:-1 , A[149], B[149], S[149]);

  wire \P149:147 , \G149:147 ;

  PijGij \149:147 (P[149], \P148:147 , G[149], \G148:147 , \P149:147 , \G149:147 );

  wire \P149:143 , \G149:143 ;

  PijGij \149:143 (\P149:147 , \P146:143 , \G149:147 , \G146:143 , \P149:143 , \G149:143 );

  wire \P149:127 , \G149:127 ;

  PijGij \149:127 (\P149:143 , \P142:127 , \G149:143 , \G142:127 , \P149:127 , \G149:127 );

  wire \G149:-1 ;

  Gij \149:-1 (\P149:127 , \G149:127 , \G126:-1 , \G149:-1 );

  Sum s150(\G149:-1 , A[150], B[150], S[150]);

  wire \P150:149 , \G150:149 ;

  PijGij \150:149 (P[150], P[149], G[150], G[149], \P150:149 , \G150:149 );

  wire \P150:147 , \G150:147 ;

  PijGij \150:147 (\P150:149 , \P148:147 , \G150:149 , \G148:147 , \P150:147 , \G150:147 );

  wire \P150:143 , \G150:143 ;

  PijGij \150:143 (\P150:147 , \P146:143 , \G150:147 , \G146:143 , \P150:143 , \G150:143 );

  wire \P150:127 , \G150:127 ;

  PijGij \150:127 (\P150:143 , \P142:127 , \G150:143 , \G142:127 , \P150:127 , \G150:127 );

  wire \G150:-1 ;

  Gij \150:-1 (\P150:127 , \G150:127 , \G126:-1 , \G150:-1 );

  Sum s151(\G150:-1 , A[151], B[151], S[151]);

  wire \P151:143 , \G151:143 ;

  PijGij \151:143 (P[151], \P150:143 , G[151], \G150:143 , \P151:143 , \G151:143 );

  wire \P151:127 , \G151:127 ;

  PijGij \151:127 (\P151:143 , \P142:127 , \G151:143 , \G142:127 , \P151:127 , \G151:127 );

  wire \G151:-1 ;

  Gij \151:-1 (\P151:127 , \G151:127 , \G126:-1 , \G151:-1 );

  Sum s152(\G151:-1 , A[152], B[152], S[152]);

  wire \P152:151 , \G152:151 ;

  PijGij \152:151 (P[152], P[151], G[152], G[151], \P152:151 , \G152:151 );

  wire \P152:143 , \G152:143 ;

  PijGij \152:143 (\P152:151 , \P150:143 , \G152:151 , \G150:143 , \P152:143 , \G152:143 );

  wire \P152:127 , \G152:127 ;

  PijGij \152:127 (\P152:143 , \P142:127 , \G152:143 , \G142:127 , \P152:127 , \G152:127 );

  wire \G152:-1 ;

  Gij \152:-1 (\P152:127 , \G152:127 , \G126:-1 , \G152:-1 );

  Sum s153(\G152:-1 , A[153], B[153], S[153]);

  wire \P153:151 , \G153:151 ;

  PijGij \153:151 (P[153], \P152:151 , G[153], \G152:151 , \P153:151 , \G153:151 );

  wire \P153:143 , \G153:143 ;

  PijGij \153:143 (\P153:151 , \P150:143 , \G153:151 , \G150:143 , \P153:143 , \G153:143 );

  wire \P153:127 , \G153:127 ;

  PijGij \153:127 (\P153:143 , \P142:127 , \G153:143 , \G142:127 , \P153:127 , \G153:127 );

  wire \G153:-1 ;

  Gij \153:-1 (\P153:127 , \G153:127 , \G126:-1 , \G153:-1 );

  Sum s154(\G153:-1 , A[154], B[154], S[154]);

  wire \P154:153 , \G154:153 ;

  PijGij \154:153 (P[154], P[153], G[154], G[153], \P154:153 , \G154:153 );

  wire \P154:151 , \G154:151 ;

  PijGij \154:151 (\P154:153 , \P152:151 , \G154:153 , \G152:151 , \P154:151 , \G154:151 );

  wire \P154:143 , \G154:143 ;

  PijGij \154:143 (\P154:151 , \P150:143 , \G154:151 , \G150:143 , \P154:143 , \G154:143 );

  wire \P154:127 , \G154:127 ;

  PijGij \154:127 (\P154:143 , \P142:127 , \G154:143 , \G142:127 , \P154:127 , \G154:127 );

  wire \G154:-1 ;

  Gij \154:-1 (\P154:127 , \G154:127 , \G126:-1 , \G154:-1 );

  Sum s155(\G154:-1 , A[155], B[155], S[155]);

  wire \P155:151 , \G155:151 ;

  PijGij \155:151 (P[155], \P154:151 , G[155], \G154:151 , \P155:151 , \G155:151 );

  wire \P155:143 , \G155:143 ;

  PijGij \155:143 (\P155:151 , \P150:143 , \G155:151 , \G150:143 , \P155:143 , \G155:143 );

  wire \P155:127 , \G155:127 ;

  PijGij \155:127 (\P155:143 , \P142:127 , \G155:143 , \G142:127 , \P155:127 , \G155:127 );

  wire \G155:-1 ;

  Gij \155:-1 (\P155:127 , \G155:127 , \G126:-1 , \G155:-1 );

  Sum s156(\G155:-1 , A[156], B[156], S[156]);

  wire \P156:155 , \G156:155 ;

  PijGij \156:155 (P[156], P[155], G[156], G[155], \P156:155 , \G156:155 );

  wire \P156:151 , \G156:151 ;

  PijGij \156:151 (\P156:155 , \P154:151 , \G156:155 , \G154:151 , \P156:151 , \G156:151 );

  wire \P156:143 , \G156:143 ;

  PijGij \156:143 (\P156:151 , \P150:143 , \G156:151 , \G150:143 , \P156:143 , \G156:143 );

  wire \P156:127 , \G156:127 ;

  PijGij \156:127 (\P156:143 , \P142:127 , \G156:143 , \G142:127 , \P156:127 , \G156:127 );

  wire \G156:-1 ;

  Gij \156:-1 (\P156:127 , \G156:127 , \G126:-1 , \G156:-1 );

  Sum s157(\G156:-1 , A[157], B[157], S[157]);

  wire \P157:155 , \G157:155 ;

  PijGij \157:155 (P[157], \P156:155 , G[157], \G156:155 , \P157:155 , \G157:155 );

  wire \P157:151 , \G157:151 ;

  PijGij \157:151 (\P157:155 , \P154:151 , \G157:155 , \G154:151 , \P157:151 , \G157:151 );

  wire \P157:143 , \G157:143 ;

  PijGij \157:143 (\P157:151 , \P150:143 , \G157:151 , \G150:143 , \P157:143 , \G157:143 );

  wire \P157:127 , \G157:127 ;

  PijGij \157:127 (\P157:143 , \P142:127 , \G157:143 , \G142:127 , \P157:127 , \G157:127 );

  wire \G157:-1 ;

  Gij \157:-1 (\P157:127 , \G157:127 , \G126:-1 , \G157:-1 );

  Sum s158(\G157:-1 , A[158], B[158], S[158]);

  wire \P158:157 , \G158:157 ;

  PijGij \158:157 (P[158], P[157], G[158], G[157], \P158:157 , \G158:157 );

  wire \P158:155 , \G158:155 ;

  PijGij \158:155 (\P158:157 , \P156:155 , \G158:157 , \G156:155 , \P158:155 , \G158:155 );

  wire \P158:151 , \G158:151 ;

  PijGij \158:151 (\P158:155 , \P154:151 , \G158:155 , \G154:151 , \P158:151 , \G158:151 );

  wire \P158:143 , \G158:143 ;

  PijGij \158:143 (\P158:151 , \P150:143 , \G158:151 , \G150:143 , \P158:143 , \G158:143 );

  wire \P158:127 , \G158:127 ;

  PijGij \158:127 (\P158:143 , \P142:127 , \G158:143 , \G142:127 , \P158:127 , \G158:127 );

  wire \G158:-1 ;

  Gij \158:-1 (\P158:127 , \G158:127 , \G126:-1 , \G158:-1 );

  Sum s159(\G158:-1 , A[159], B[159], S[159]);

  wire \P159:127 , \G159:127 ;

  PijGij \159:127 (P[159], \P158:127 , G[159], \G158:127 , \P159:127 , \G159:127 );

  wire \G159:-1 ;

  Gij \159:-1 (\P159:127 , \G159:127 , \G126:-1 , \G159:-1 );

  Sum s160(\G159:-1 , A[160], B[160], S[160]);

  wire \P160:159 , \G160:159 ;

  PijGij \160:159 (P[160], P[159], G[160], G[159], \P160:159 , \G160:159 );

  wire \P160:127 , \G160:127 ;

  PijGij \160:127 (\P160:159 , \P158:127 , \G160:159 , \G158:127 , \P160:127 , \G160:127 );

  wire \G160:-1 ;

  Gij \160:-1 (\P160:127 , \G160:127 , \G126:-1 , \G160:-1 );

  Sum s161(\G160:-1 , A[161], B[161], S[161]);

  wire \P161:159 , \G161:159 ;

  PijGij \161:159 (P[161], \P160:159 , G[161], \G160:159 , \P161:159 , \G161:159 );

  wire \P161:127 , \G161:127 ;

  PijGij \161:127 (\P161:159 , \P158:127 , \G161:159 , \G158:127 , \P161:127 , \G161:127 );

  wire \G161:-1 ;

  Gij \161:-1 (\P161:127 , \G161:127 , \G126:-1 , \G161:-1 );

  Sum s162(\G161:-1 , A[162], B[162], S[162]);

  wire \P162:161 , \G162:161 ;

  PijGij \162:161 (P[162], P[161], G[162], G[161], \P162:161 , \G162:161 );

  wire \P162:159 , \G162:159 ;

  PijGij \162:159 (\P162:161 , \P160:159 , \G162:161 , \G160:159 , \P162:159 , \G162:159 );

  wire \P162:127 , \G162:127 ;

  PijGij \162:127 (\P162:159 , \P158:127 , \G162:159 , \G158:127 , \P162:127 , \G162:127 );

  wire \G162:-1 ;

  Gij \162:-1 (\P162:127 , \G162:127 , \G126:-1 , \G162:-1 );

  Sum s163(\G162:-1 , A[163], B[163], S[163]);

  wire \P163:159 , \G163:159 ;

  PijGij \163:159 (P[163], \P162:159 , G[163], \G162:159 , \P163:159 , \G163:159 );

  wire \P163:127 , \G163:127 ;

  PijGij \163:127 (\P163:159 , \P158:127 , \G163:159 , \G158:127 , \P163:127 , \G163:127 );

  wire \G163:-1 ;

  Gij \163:-1 (\P163:127 , \G163:127 , \G126:-1 , \G163:-1 );

  Sum s164(\G163:-1 , A[164], B[164], S[164]);

  wire \P164:163 , \G164:163 ;

  PijGij \164:163 (P[164], P[163], G[164], G[163], \P164:163 , \G164:163 );

  wire \P164:159 , \G164:159 ;

  PijGij \164:159 (\P164:163 , \P162:159 , \G164:163 , \G162:159 , \P164:159 , \G164:159 );

  wire \P164:127 , \G164:127 ;

  PijGij \164:127 (\P164:159 , \P158:127 , \G164:159 , \G158:127 , \P164:127 , \G164:127 );

  wire \G164:-1 ;

  Gij \164:-1 (\P164:127 , \G164:127 , \G126:-1 , \G164:-1 );

  Sum s165(\G164:-1 , A[165], B[165], S[165]);

  wire \P165:163 , \G165:163 ;

  PijGij \165:163 (P[165], \P164:163 , G[165], \G164:163 , \P165:163 , \G165:163 );

  wire \P165:159 , \G165:159 ;

  PijGij \165:159 (\P165:163 , \P162:159 , \G165:163 , \G162:159 , \P165:159 , \G165:159 );

  wire \P165:127 , \G165:127 ;

  PijGij \165:127 (\P165:159 , \P158:127 , \G165:159 , \G158:127 , \P165:127 , \G165:127 );

  wire \G165:-1 ;

  Gij \165:-1 (\P165:127 , \G165:127 , \G126:-1 , \G165:-1 );

  Sum s166(\G165:-1 , A[166], B[166], S[166]);

  wire \P166:165 , \G166:165 ;

  PijGij \166:165 (P[166], P[165], G[166], G[165], \P166:165 , \G166:165 );

  wire \P166:163 , \G166:163 ;

  PijGij \166:163 (\P166:165 , \P164:163 , \G166:165 , \G164:163 , \P166:163 , \G166:163 );

  wire \P166:159 , \G166:159 ;

  PijGij \166:159 (\P166:163 , \P162:159 , \G166:163 , \G162:159 , \P166:159 , \G166:159 );

  wire \P166:127 , \G166:127 ;

  PijGij \166:127 (\P166:159 , \P158:127 , \G166:159 , \G158:127 , \P166:127 , \G166:127 );

  wire \G166:-1 ;

  Gij \166:-1 (\P166:127 , \G166:127 , \G126:-1 , \G166:-1 );

  Sum s167(\G166:-1 , A[167], B[167], S[167]);

  wire \P167:159 , \G167:159 ;

  PijGij \167:159 (P[167], \P166:159 , G[167], \G166:159 , \P167:159 , \G167:159 );

  wire \P167:127 , \G167:127 ;

  PijGij \167:127 (\P167:159 , \P158:127 , \G167:159 , \G158:127 , \P167:127 , \G167:127 );

  wire \G167:-1 ;

  Gij \167:-1 (\P167:127 , \G167:127 , \G126:-1 , \G167:-1 );

  Sum s168(\G167:-1 , A[168], B[168], S[168]);

  wire \P168:167 , \G168:167 ;

  PijGij \168:167 (P[168], P[167], G[168], G[167], \P168:167 , \G168:167 );

  wire \P168:159 , \G168:159 ;

  PijGij \168:159 (\P168:167 , \P166:159 , \G168:167 , \G166:159 , \P168:159 , \G168:159 );

  wire \P168:127 , \G168:127 ;

  PijGij \168:127 (\P168:159 , \P158:127 , \G168:159 , \G158:127 , \P168:127 , \G168:127 );

  wire \G168:-1 ;

  Gij \168:-1 (\P168:127 , \G168:127 , \G126:-1 , \G168:-1 );

  Sum s169(\G168:-1 , A[169], B[169], S[169]);

  wire \P169:167 , \G169:167 ;

  PijGij \169:167 (P[169], \P168:167 , G[169], \G168:167 , \P169:167 , \G169:167 );

  wire \P169:159 , \G169:159 ;

  PijGij \169:159 (\P169:167 , \P166:159 , \G169:167 , \G166:159 , \P169:159 , \G169:159 );

  wire \P169:127 , \G169:127 ;

  PijGij \169:127 (\P169:159 , \P158:127 , \G169:159 , \G158:127 , \P169:127 , \G169:127 );

  wire \G169:-1 ;

  Gij \169:-1 (\P169:127 , \G169:127 , \G126:-1 , \G169:-1 );

  Sum s170(\G169:-1 , A[170], B[170], S[170]);

  wire \P170:169 , \G170:169 ;

  PijGij \170:169 (P[170], P[169], G[170], G[169], \P170:169 , \G170:169 );

  wire \P170:167 , \G170:167 ;

  PijGij \170:167 (\P170:169 , \P168:167 , \G170:169 , \G168:167 , \P170:167 , \G170:167 );

  wire \P170:159 , \G170:159 ;

  PijGij \170:159 (\P170:167 , \P166:159 , \G170:167 , \G166:159 , \P170:159 , \G170:159 );

  wire \P170:127 , \G170:127 ;

  PijGij \170:127 (\P170:159 , \P158:127 , \G170:159 , \G158:127 , \P170:127 , \G170:127 );

  wire \G170:-1 ;

  Gij \170:-1 (\P170:127 , \G170:127 , \G126:-1 , \G170:-1 );

  Sum s171(\G170:-1 , A[171], B[171], S[171]);

  wire \P171:167 , \G171:167 ;

  PijGij \171:167 (P[171], \P170:167 , G[171], \G170:167 , \P171:167 , \G171:167 );

  wire \P171:159 , \G171:159 ;

  PijGij \171:159 (\P171:167 , \P166:159 , \G171:167 , \G166:159 , \P171:159 , \G171:159 );

  wire \P171:127 , \G171:127 ;

  PijGij \171:127 (\P171:159 , \P158:127 , \G171:159 , \G158:127 , \P171:127 , \G171:127 );

  wire \G171:-1 ;

  Gij \171:-1 (\P171:127 , \G171:127 , \G126:-1 , \G171:-1 );

  Sum s172(\G171:-1 , A[172], B[172], S[172]);

  wire \P172:171 , \G172:171 ;

  PijGij \172:171 (P[172], P[171], G[172], G[171], \P172:171 , \G172:171 );

  wire \P172:167 , \G172:167 ;

  PijGij \172:167 (\P172:171 , \P170:167 , \G172:171 , \G170:167 , \P172:167 , \G172:167 );

  wire \P172:159 , \G172:159 ;

  PijGij \172:159 (\P172:167 , \P166:159 , \G172:167 , \G166:159 , \P172:159 , \G172:159 );

  wire \P172:127 , \G172:127 ;

  PijGij \172:127 (\P172:159 , \P158:127 , \G172:159 , \G158:127 , \P172:127 , \G172:127 );

  wire \G172:-1 ;

  Gij \172:-1 (\P172:127 , \G172:127 , \G126:-1 , \G172:-1 );

  Sum s173(\G172:-1 , A[173], B[173], S[173]);

  wire \P173:171 , \G173:171 ;

  PijGij \173:171 (P[173], \P172:171 , G[173], \G172:171 , \P173:171 , \G173:171 );

  wire \P173:167 , \G173:167 ;

  PijGij \173:167 (\P173:171 , \P170:167 , \G173:171 , \G170:167 , \P173:167 , \G173:167 );

  wire \P173:159 , \G173:159 ;

  PijGij \173:159 (\P173:167 , \P166:159 , \G173:167 , \G166:159 , \P173:159 , \G173:159 );

  wire \P173:127 , \G173:127 ;

  PijGij \173:127 (\P173:159 , \P158:127 , \G173:159 , \G158:127 , \P173:127 , \G173:127 );

  wire \G173:-1 ;

  Gij \173:-1 (\P173:127 , \G173:127 , \G126:-1 , \G173:-1 );

  Sum s174(\G173:-1 , A[174], B[174], S[174]);

  wire \P174:173 , \G174:173 ;

  PijGij \174:173 (P[174], P[173], G[174], G[173], \P174:173 , \G174:173 );

  wire \P174:171 , \G174:171 ;

  PijGij \174:171 (\P174:173 , \P172:171 , \G174:173 , \G172:171 , \P174:171 , \G174:171 );

  wire \P174:167 , \G174:167 ;

  PijGij \174:167 (\P174:171 , \P170:167 , \G174:171 , \G170:167 , \P174:167 , \G174:167 );

  wire \P174:159 , \G174:159 ;

  PijGij \174:159 (\P174:167 , \P166:159 , \G174:167 , \G166:159 , \P174:159 , \G174:159 );

  wire \P174:127 , \G174:127 ;

  PijGij \174:127 (\P174:159 , \P158:127 , \G174:159 , \G158:127 , \P174:127 , \G174:127 );

  wire \G174:-1 ;

  Gij \174:-1 (\P174:127 , \G174:127 , \G126:-1 , \G174:-1 );

  Sum s175(\G174:-1 , A[175], B[175], S[175]);

  wire \P175:159 , \G175:159 ;

  PijGij \175:159 (P[175], \P174:159 , G[175], \G174:159 , \P175:159 , \G175:159 );

  wire \P175:127 , \G175:127 ;

  PijGij \175:127 (\P175:159 , \P158:127 , \G175:159 , \G158:127 , \P175:127 , \G175:127 );

  wire \G175:-1 ;

  Gij \175:-1 (\P175:127 , \G175:127 , \G126:-1 , \G175:-1 );

  Sum s176(\G175:-1 , A[176], B[176], S[176]);

  wire \P176:175 , \G176:175 ;

  PijGij \176:175 (P[176], P[175], G[176], G[175], \P176:175 , \G176:175 );

  wire \P176:159 , \G176:159 ;

  PijGij \176:159 (\P176:175 , \P174:159 , \G176:175 , \G174:159 , \P176:159 , \G176:159 );

  wire \P176:127 , \G176:127 ;

  PijGij \176:127 (\P176:159 , \P158:127 , \G176:159 , \G158:127 , \P176:127 , \G176:127 );

  wire \G176:-1 ;

  Gij \176:-1 (\P176:127 , \G176:127 , \G126:-1 , \G176:-1 );

  Sum s177(\G176:-1 , A[177], B[177], S[177]);

  wire \P177:175 , \G177:175 ;

  PijGij \177:175 (P[177], \P176:175 , G[177], \G176:175 , \P177:175 , \G177:175 );

  wire \P177:159 , \G177:159 ;

  PijGij \177:159 (\P177:175 , \P174:159 , \G177:175 , \G174:159 , \P177:159 , \G177:159 );

  wire \P177:127 , \G177:127 ;

  PijGij \177:127 (\P177:159 , \P158:127 , \G177:159 , \G158:127 , \P177:127 , \G177:127 );

  wire \G177:-1 ;

  Gij \177:-1 (\P177:127 , \G177:127 , \G126:-1 , \G177:-1 );

  Sum s178(\G177:-1 , A[178], B[178], S[178]);

  wire \P178:177 , \G178:177 ;

  PijGij \178:177 (P[178], P[177], G[178], G[177], \P178:177 , \G178:177 );

  wire \P178:175 , \G178:175 ;

  PijGij \178:175 (\P178:177 , \P176:175 , \G178:177 , \G176:175 , \P178:175 , \G178:175 );

  wire \P178:159 , \G178:159 ;

  PijGij \178:159 (\P178:175 , \P174:159 , \G178:175 , \G174:159 , \P178:159 , \G178:159 );

  wire \P178:127 , \G178:127 ;

  PijGij \178:127 (\P178:159 , \P158:127 , \G178:159 , \G158:127 , \P178:127 , \G178:127 );

  wire \G178:-1 ;

  Gij \178:-1 (\P178:127 , \G178:127 , \G126:-1 , \G178:-1 );

  Sum s179(\G178:-1 , A[179], B[179], S[179]);

  wire \P179:175 , \G179:175 ;

  PijGij \179:175 (P[179], \P178:175 , G[179], \G178:175 , \P179:175 , \G179:175 );

  wire \P179:159 , \G179:159 ;

  PijGij \179:159 (\P179:175 , \P174:159 , \G179:175 , \G174:159 , \P179:159 , \G179:159 );

  wire \P179:127 , \G179:127 ;

  PijGij \179:127 (\P179:159 , \P158:127 , \G179:159 , \G158:127 , \P179:127 , \G179:127 );

  wire \G179:-1 ;

  Gij \179:-1 (\P179:127 , \G179:127 , \G126:-1 , \G179:-1 );

  Sum s180(\G179:-1 , A[180], B[180], S[180]);

  wire \P180:179 , \G180:179 ;

  PijGij \180:179 (P[180], P[179], G[180], G[179], \P180:179 , \G180:179 );

  wire \P180:175 , \G180:175 ;

  PijGij \180:175 (\P180:179 , \P178:175 , \G180:179 , \G178:175 , \P180:175 , \G180:175 );

  wire \P180:159 , \G180:159 ;

  PijGij \180:159 (\P180:175 , \P174:159 , \G180:175 , \G174:159 , \P180:159 , \G180:159 );

  wire \P180:127 , \G180:127 ;

  PijGij \180:127 (\P180:159 , \P158:127 , \G180:159 , \G158:127 , \P180:127 , \G180:127 );

  wire \G180:-1 ;

  Gij \180:-1 (\P180:127 , \G180:127 , \G126:-1 , \G180:-1 );

  Sum s181(\G180:-1 , A[181], B[181], S[181]);

  wire \P181:179 , \G181:179 ;

  PijGij \181:179 (P[181], \P180:179 , G[181], \G180:179 , \P181:179 , \G181:179 );

  wire \P181:175 , \G181:175 ;

  PijGij \181:175 (\P181:179 , \P178:175 , \G181:179 , \G178:175 , \P181:175 , \G181:175 );

  wire \P181:159 , \G181:159 ;

  PijGij \181:159 (\P181:175 , \P174:159 , \G181:175 , \G174:159 , \P181:159 , \G181:159 );

  wire \P181:127 , \G181:127 ;

  PijGij \181:127 (\P181:159 , \P158:127 , \G181:159 , \G158:127 , \P181:127 , \G181:127 );

  wire \G181:-1 ;

  Gij \181:-1 (\P181:127 , \G181:127 , \G126:-1 , \G181:-1 );

  Sum s182(\G181:-1 , A[182], B[182], S[182]);

  wire \P182:181 , \G182:181 ;

  PijGij \182:181 (P[182], P[181], G[182], G[181], \P182:181 , \G182:181 );

  wire \P182:179 , \G182:179 ;

  PijGij \182:179 (\P182:181 , \P180:179 , \G182:181 , \G180:179 , \P182:179 , \G182:179 );

  wire \P182:175 , \G182:175 ;

  PijGij \182:175 (\P182:179 , \P178:175 , \G182:179 , \G178:175 , \P182:175 , \G182:175 );

  wire \P182:159 , \G182:159 ;

  PijGij \182:159 (\P182:175 , \P174:159 , \G182:175 , \G174:159 , \P182:159 , \G182:159 );

  wire \P182:127 , \G182:127 ;

  PijGij \182:127 (\P182:159 , \P158:127 , \G182:159 , \G158:127 , \P182:127 , \G182:127 );

  wire \G182:-1 ;

  Gij \182:-1 (\P182:127 , \G182:127 , \G126:-1 , \G182:-1 );

  Sum s183(\G182:-1 , A[183], B[183], S[183]);

  wire \P183:175 , \G183:175 ;

  PijGij \183:175 (P[183], \P182:175 , G[183], \G182:175 , \P183:175 , \G183:175 );

  wire \P183:159 , \G183:159 ;

  PijGij \183:159 (\P183:175 , \P174:159 , \G183:175 , \G174:159 , \P183:159 , \G183:159 );

  wire \P183:127 , \G183:127 ;

  PijGij \183:127 (\P183:159 , \P158:127 , \G183:159 , \G158:127 , \P183:127 , \G183:127 );

  wire \G183:-1 ;

  Gij \183:-1 (\P183:127 , \G183:127 , \G126:-1 , \G183:-1 );

  Sum s184(\G183:-1 , A[184], B[184], S[184]);

  wire \P184:183 , \G184:183 ;

  PijGij \184:183 (P[184], P[183], G[184], G[183], \P184:183 , \G184:183 );

  wire \P184:175 , \G184:175 ;

  PijGij \184:175 (\P184:183 , \P182:175 , \G184:183 , \G182:175 , \P184:175 , \G184:175 );

  wire \P184:159 , \G184:159 ;

  PijGij \184:159 (\P184:175 , \P174:159 , \G184:175 , \G174:159 , \P184:159 , \G184:159 );

  wire \P184:127 , \G184:127 ;

  PijGij \184:127 (\P184:159 , \P158:127 , \G184:159 , \G158:127 , \P184:127 , \G184:127 );

  wire \G184:-1 ;

  Gij \184:-1 (\P184:127 , \G184:127 , \G126:-1 , \G184:-1 );

  Sum s185(\G184:-1 , A[185], B[185], S[185]);

  wire \P185:183 , \G185:183 ;

  PijGij \185:183 (P[185], \P184:183 , G[185], \G184:183 , \P185:183 , \G185:183 );

  wire \P185:175 , \G185:175 ;

  PijGij \185:175 (\P185:183 , \P182:175 , \G185:183 , \G182:175 , \P185:175 , \G185:175 );

  wire \P185:159 , \G185:159 ;

  PijGij \185:159 (\P185:175 , \P174:159 , \G185:175 , \G174:159 , \P185:159 , \G185:159 );

  wire \P185:127 , \G185:127 ;

  PijGij \185:127 (\P185:159 , \P158:127 , \G185:159 , \G158:127 , \P185:127 , \G185:127 );

  wire \G185:-1 ;

  Gij \185:-1 (\P185:127 , \G185:127 , \G126:-1 , \G185:-1 );

  Sum s186(\G185:-1 , A[186], B[186], S[186]);

  wire \P186:185 , \G186:185 ;

  PijGij \186:185 (P[186], P[185], G[186], G[185], \P186:185 , \G186:185 );

  wire \P186:183 , \G186:183 ;

  PijGij \186:183 (\P186:185 , \P184:183 , \G186:185 , \G184:183 , \P186:183 , \G186:183 );

  wire \P186:175 , \G186:175 ;

  PijGij \186:175 (\P186:183 , \P182:175 , \G186:183 , \G182:175 , \P186:175 , \G186:175 );

  wire \P186:159 , \G186:159 ;

  PijGij \186:159 (\P186:175 , \P174:159 , \G186:175 , \G174:159 , \P186:159 , \G186:159 );

  wire \P186:127 , \G186:127 ;

  PijGij \186:127 (\P186:159 , \P158:127 , \G186:159 , \G158:127 , \P186:127 , \G186:127 );

  wire \G186:-1 ;

  Gij \186:-1 (\P186:127 , \G186:127 , \G126:-1 , \G186:-1 );

  Sum s187(\G186:-1 , A[187], B[187], S[187]);

  wire \P187:183 , \G187:183 ;

  PijGij \187:183 (P[187], \P186:183 , G[187], \G186:183 , \P187:183 , \G187:183 );

  wire \P187:175 , \G187:175 ;

  PijGij \187:175 (\P187:183 , \P182:175 , \G187:183 , \G182:175 , \P187:175 , \G187:175 );

  wire \P187:159 , \G187:159 ;

  PijGij \187:159 (\P187:175 , \P174:159 , \G187:175 , \G174:159 , \P187:159 , \G187:159 );

  wire \P187:127 , \G187:127 ;

  PijGij \187:127 (\P187:159 , \P158:127 , \G187:159 , \G158:127 , \P187:127 , \G187:127 );

  wire \G187:-1 ;

  Gij \187:-1 (\P187:127 , \G187:127 , \G126:-1 , \G187:-1 );

  Sum s188(\G187:-1 , A[188], B[188], S[188]);

  wire \P188:187 , \G188:187 ;

  PijGij \188:187 (P[188], P[187], G[188], G[187], \P188:187 , \G188:187 );

  wire \P188:183 , \G188:183 ;

  PijGij \188:183 (\P188:187 , \P186:183 , \G188:187 , \G186:183 , \P188:183 , \G188:183 );

  wire \P188:175 , \G188:175 ;

  PijGij \188:175 (\P188:183 , \P182:175 , \G188:183 , \G182:175 , \P188:175 , \G188:175 );

  wire \P188:159 , \G188:159 ;

  PijGij \188:159 (\P188:175 , \P174:159 , \G188:175 , \G174:159 , \P188:159 , \G188:159 );

  wire \P188:127 , \G188:127 ;

  PijGij \188:127 (\P188:159 , \P158:127 , \G188:159 , \G158:127 , \P188:127 , \G188:127 );

  wire \G188:-1 ;

  Gij \188:-1 (\P188:127 , \G188:127 , \G126:-1 , \G188:-1 );

  Sum s189(\G188:-1 , A[189], B[189], S[189]);

  wire \P189:187 , \G189:187 ;

  PijGij \189:187 (P[189], \P188:187 , G[189], \G188:187 , \P189:187 , \G189:187 );

  wire \P189:183 , \G189:183 ;

  PijGij \189:183 (\P189:187 , \P186:183 , \G189:187 , \G186:183 , \P189:183 , \G189:183 );

  wire \P189:175 , \G189:175 ;

  PijGij \189:175 (\P189:183 , \P182:175 , \G189:183 , \G182:175 , \P189:175 , \G189:175 );

  wire \P189:159 , \G189:159 ;

  PijGij \189:159 (\P189:175 , \P174:159 , \G189:175 , \G174:159 , \P189:159 , \G189:159 );

  wire \P189:127 , \G189:127 ;

  PijGij \189:127 (\P189:159 , \P158:127 , \G189:159 , \G158:127 , \P189:127 , \G189:127 );

  wire \G189:-1 ;

  Gij \189:-1 (\P189:127 , \G189:127 , \G126:-1 , \G189:-1 );

  Sum s190(\G189:-1 , A[190], B[190], S[190]);

  wire \P190:189 , \G190:189 ;

  PijGij \190:189 (P[190], P[189], G[190], G[189], \P190:189 , \G190:189 );

  wire \P190:187 , \G190:187 ;

  PijGij \190:187 (\P190:189 , \P188:187 , \G190:189 , \G188:187 , \P190:187 , \G190:187 );

  wire \P190:183 , \G190:183 ;

  PijGij \190:183 (\P190:187 , \P186:183 , \G190:187 , \G186:183 , \P190:183 , \G190:183 );

  wire \P190:175 , \G190:175 ;

  PijGij \190:175 (\P190:183 , \P182:175 , \G190:183 , \G182:175 , \P190:175 , \G190:175 );

  wire \P190:159 , \G190:159 ;

  PijGij \190:159 (\P190:175 , \P174:159 , \G190:175 , \G174:159 , \P190:159 , \G190:159 );

  wire \P190:127 , \G190:127 ;

  PijGij \190:127 (\P190:159 , \P158:127 , \G190:159 , \G158:127 , \P190:127 , \G190:127 );

  wire \G190:-1 ;

  Gij \190:-1 (\P190:127 , \G190:127 , \G126:-1 , \G190:-1 );

  Sum s191(\G190:-1 , A[191], B[191], S[191]);

  wire \P191:127 , \G191:127 ;

  PijGij \191:127 (P[191], \P190:127 , G[191], \G190:127 , \P191:127 , \G191:127 );

  wire \G191:-1 ;

  Gij \191:-1 (\P191:127 , \G191:127 , \G126:-1 , \G191:-1 );

  Sum s192(\G191:-1 , A[192], B[192], S[192]);

  wire \P192:191 , \G192:191 ;

  PijGij \192:191 (P[192], P[191], G[192], G[191], \P192:191 , \G192:191 );

  wire \P192:127 , \G192:127 ;

  PijGij \192:127 (\P192:191 , \P190:127 , \G192:191 , \G190:127 , \P192:127 , \G192:127 );

  wire \G192:-1 ;

  Gij \192:-1 (\P192:127 , \G192:127 , \G126:-1 , \G192:-1 );

  Sum s193(\G192:-1 , A[193], B[193], S[193]);

  wire \P193:191 , \G193:191 ;

  PijGij \193:191 (P[193], \P192:191 , G[193], \G192:191 , \P193:191 , \G193:191 );

  wire \P193:127 , \G193:127 ;

  PijGij \193:127 (\P193:191 , \P190:127 , \G193:191 , \G190:127 , \P193:127 , \G193:127 );

  wire \G193:-1 ;

  Gij \193:-1 (\P193:127 , \G193:127 , \G126:-1 , \G193:-1 );

  Sum s194(\G193:-1 , A[194], B[194], S[194]);

  wire \P194:193 , \G194:193 ;

  PijGij \194:193 (P[194], P[193], G[194], G[193], \P194:193 , \G194:193 );

  wire \P194:191 , \G194:191 ;

  PijGij \194:191 (\P194:193 , \P192:191 , \G194:193 , \G192:191 , \P194:191 , \G194:191 );

  wire \P194:127 , \G194:127 ;

  PijGij \194:127 (\P194:191 , \P190:127 , \G194:191 , \G190:127 , \P194:127 , \G194:127 );

  wire \G194:-1 ;

  Gij \194:-1 (\P194:127 , \G194:127 , \G126:-1 , \G194:-1 );

  Sum s195(\G194:-1 , A[195], B[195], S[195]);

  wire \P195:191 , \G195:191 ;

  PijGij \195:191 (P[195], \P194:191 , G[195], \G194:191 , \P195:191 , \G195:191 );

  wire \P195:127 , \G195:127 ;

  PijGij \195:127 (\P195:191 , \P190:127 , \G195:191 , \G190:127 , \P195:127 , \G195:127 );

  wire \G195:-1 ;

  Gij \195:-1 (\P195:127 , \G195:127 , \G126:-1 , \G195:-1 );

  Sum s196(\G195:-1 , A[196], B[196], S[196]);

  wire \P196:195 , \G196:195 ;

  PijGij \196:195 (P[196], P[195], G[196], G[195], \P196:195 , \G196:195 );

  wire \P196:191 , \G196:191 ;

  PijGij \196:191 (\P196:195 , \P194:191 , \G196:195 , \G194:191 , \P196:191 , \G196:191 );

  wire \P196:127 , \G196:127 ;

  PijGij \196:127 (\P196:191 , \P190:127 , \G196:191 , \G190:127 , \P196:127 , \G196:127 );

  wire \G196:-1 ;

  Gij \196:-1 (\P196:127 , \G196:127 , \G126:-1 , \G196:-1 );

  Sum s197(\G196:-1 , A[197], B[197], S[197]);

  wire \P197:195 , \G197:195 ;

  PijGij \197:195 (P[197], \P196:195 , G[197], \G196:195 , \P197:195 , \G197:195 );

  wire \P197:191 , \G197:191 ;

  PijGij \197:191 (\P197:195 , \P194:191 , \G197:195 , \G194:191 , \P197:191 , \G197:191 );

  wire \P197:127 , \G197:127 ;

  PijGij \197:127 (\P197:191 , \P190:127 , \G197:191 , \G190:127 , \P197:127 , \G197:127 );

  wire \G197:-1 ;

  Gij \197:-1 (\P197:127 , \G197:127 , \G126:-1 , \G197:-1 );

  Sum s198(\G197:-1 , A[198], B[198], S[198]);

  wire \P198:197 , \G198:197 ;

  PijGij \198:197 (P[198], P[197], G[198], G[197], \P198:197 , \G198:197 );

  wire \P198:195 , \G198:195 ;

  PijGij \198:195 (\P198:197 , \P196:195 , \G198:197 , \G196:195 , \P198:195 , \G198:195 );

  wire \P198:191 , \G198:191 ;

  PijGij \198:191 (\P198:195 , \P194:191 , \G198:195 , \G194:191 , \P198:191 , \G198:191 );

  wire \P198:127 , \G198:127 ;

  PijGij \198:127 (\P198:191 , \P190:127 , \G198:191 , \G190:127 , \P198:127 , \G198:127 );

  wire \G198:-1 ;

  Gij \198:-1 (\P198:127 , \G198:127 , \G126:-1 , \G198:-1 );

  Sum s199(\G198:-1 , A[199], B[199], S[199]);

  wire \P199:191 , \G199:191 ;

  PijGij \199:191 (P[199], \P198:191 , G[199], \G198:191 , \P199:191 , \G199:191 );

  wire \P199:127 , \G199:127 ;

  PijGij \199:127 (\P199:191 , \P190:127 , \G199:191 , \G190:127 , \P199:127 , \G199:127 );

  wire \G199:-1 ;

  Gij \199:-1 (\P199:127 , \G199:127 , \G126:-1 , \G199:-1 );

  Sum s200(\G199:-1 , A[200], B[200], S[200]);

  wire \P200:199 , \G200:199 ;

  PijGij \200:199 (P[200], P[199], G[200], G[199], \P200:199 , \G200:199 );

  wire \P200:191 , \G200:191 ;

  PijGij \200:191 (\P200:199 , \P198:191 , \G200:199 , \G198:191 , \P200:191 , \G200:191 );

  wire \P200:127 , \G200:127 ;

  PijGij \200:127 (\P200:191 , \P190:127 , \G200:191 , \G190:127 , \P200:127 , \G200:127 );

  wire \G200:-1 ;

  Gij \200:-1 (\P200:127 , \G200:127 , \G126:-1 , \G200:-1 );

  Sum s201(\G200:-1 , A[201], B[201], S[201]);

  wire \P201:199 , \G201:199 ;

  PijGij \201:199 (P[201], \P200:199 , G[201], \G200:199 , \P201:199 , \G201:199 );

  wire \P201:191 , \G201:191 ;

  PijGij \201:191 (\P201:199 , \P198:191 , \G201:199 , \G198:191 , \P201:191 , \G201:191 );

  wire \P201:127 , \G201:127 ;

  PijGij \201:127 (\P201:191 , \P190:127 , \G201:191 , \G190:127 , \P201:127 , \G201:127 );

  wire \G201:-1 ;

  Gij \201:-1 (\P201:127 , \G201:127 , \G126:-1 , \G201:-1 );

  Sum s202(\G201:-1 , A[202], B[202], S[202]);

  wire \P202:201 , \G202:201 ;

  PijGij \202:201 (P[202], P[201], G[202], G[201], \P202:201 , \G202:201 );

  wire \P202:199 , \G202:199 ;

  PijGij \202:199 (\P202:201 , \P200:199 , \G202:201 , \G200:199 , \P202:199 , \G202:199 );

  wire \P202:191 , \G202:191 ;

  PijGij \202:191 (\P202:199 , \P198:191 , \G202:199 , \G198:191 , \P202:191 , \G202:191 );

  wire \P202:127 , \G202:127 ;

  PijGij \202:127 (\P202:191 , \P190:127 , \G202:191 , \G190:127 , \P202:127 , \G202:127 );

  wire \G202:-1 ;

  Gij \202:-1 (\P202:127 , \G202:127 , \G126:-1 , \G202:-1 );

  Sum s203(\G202:-1 , A[203], B[203], S[203]);

  wire \P203:199 , \G203:199 ;

  PijGij \203:199 (P[203], \P202:199 , G[203], \G202:199 , \P203:199 , \G203:199 );

  wire \P203:191 , \G203:191 ;

  PijGij \203:191 (\P203:199 , \P198:191 , \G203:199 , \G198:191 , \P203:191 , \G203:191 );

  wire \P203:127 , \G203:127 ;

  PijGij \203:127 (\P203:191 , \P190:127 , \G203:191 , \G190:127 , \P203:127 , \G203:127 );

  wire \G203:-1 ;

  Gij \203:-1 (\P203:127 , \G203:127 , \G126:-1 , \G203:-1 );

  Sum s204(\G203:-1 , A[204], B[204], S[204]);

  wire \P204:203 , \G204:203 ;

  PijGij \204:203 (P[204], P[203], G[204], G[203], \P204:203 , \G204:203 );

  wire \P204:199 , \G204:199 ;

  PijGij \204:199 (\P204:203 , \P202:199 , \G204:203 , \G202:199 , \P204:199 , \G204:199 );

  wire \P204:191 , \G204:191 ;

  PijGij \204:191 (\P204:199 , \P198:191 , \G204:199 , \G198:191 , \P204:191 , \G204:191 );

  wire \P204:127 , \G204:127 ;

  PijGij \204:127 (\P204:191 , \P190:127 , \G204:191 , \G190:127 , \P204:127 , \G204:127 );

  wire \G204:-1 ;

  Gij \204:-1 (\P204:127 , \G204:127 , \G126:-1 , \G204:-1 );

  Sum s205(\G204:-1 , A[205], B[205], S[205]);

  wire \P205:203 , \G205:203 ;

  PijGij \205:203 (P[205], \P204:203 , G[205], \G204:203 , \P205:203 , \G205:203 );

  wire \P205:199 , \G205:199 ;

  PijGij \205:199 (\P205:203 , \P202:199 , \G205:203 , \G202:199 , \P205:199 , \G205:199 );

  wire \P205:191 , \G205:191 ;

  PijGij \205:191 (\P205:199 , \P198:191 , \G205:199 , \G198:191 , \P205:191 , \G205:191 );

  wire \P205:127 , \G205:127 ;

  PijGij \205:127 (\P205:191 , \P190:127 , \G205:191 , \G190:127 , \P205:127 , \G205:127 );

  wire \G205:-1 ;

  Gij \205:-1 (\P205:127 , \G205:127 , \G126:-1 , \G205:-1 );

  Sum s206(\G205:-1 , A[206], B[206], S[206]);

  wire \P206:205 , \G206:205 ;

  PijGij \206:205 (P[206], P[205], G[206], G[205], \P206:205 , \G206:205 );

  wire \P206:203 , \G206:203 ;

  PijGij \206:203 (\P206:205 , \P204:203 , \G206:205 , \G204:203 , \P206:203 , \G206:203 );

  wire \P206:199 , \G206:199 ;

  PijGij \206:199 (\P206:203 , \P202:199 , \G206:203 , \G202:199 , \P206:199 , \G206:199 );

  wire \P206:191 , \G206:191 ;

  PijGij \206:191 (\P206:199 , \P198:191 , \G206:199 , \G198:191 , \P206:191 , \G206:191 );

  wire \P206:127 , \G206:127 ;

  PijGij \206:127 (\P206:191 , \P190:127 , \G206:191 , \G190:127 , \P206:127 , \G206:127 );

  wire \G206:-1 ;

  Gij \206:-1 (\P206:127 , \G206:127 , \G126:-1 , \G206:-1 );

  Sum s207(\G206:-1 , A[207], B[207], S[207]);

  wire \P207:191 , \G207:191 ;

  PijGij \207:191 (P[207], \P206:191 , G[207], \G206:191 , \P207:191 , \G207:191 );

  wire \P207:127 , \G207:127 ;

  PijGij \207:127 (\P207:191 , \P190:127 , \G207:191 , \G190:127 , \P207:127 , \G207:127 );

  wire \G207:-1 ;

  Gij \207:-1 (\P207:127 , \G207:127 , \G126:-1 , \G207:-1 );

  Sum s208(\G207:-1 , A[208], B[208], S[208]);

  wire \P208:207 , \G208:207 ;

  PijGij \208:207 (P[208], P[207], G[208], G[207], \P208:207 , \G208:207 );

  wire \P208:191 , \G208:191 ;

  PijGij \208:191 (\P208:207 , \P206:191 , \G208:207 , \G206:191 , \P208:191 , \G208:191 );

  wire \P208:127 , \G208:127 ;

  PijGij \208:127 (\P208:191 , \P190:127 , \G208:191 , \G190:127 , \P208:127 , \G208:127 );

  wire \G208:-1 ;

  Gij \208:-1 (\P208:127 , \G208:127 , \G126:-1 , \G208:-1 );

  Sum s209(\G208:-1 , A[209], B[209], S[209]);

  wire \P209:207 , \G209:207 ;

  PijGij \209:207 (P[209], \P208:207 , G[209], \G208:207 , \P209:207 , \G209:207 );

  wire \P209:191 , \G209:191 ;

  PijGij \209:191 (\P209:207 , \P206:191 , \G209:207 , \G206:191 , \P209:191 , \G209:191 );

  wire \P209:127 , \G209:127 ;

  PijGij \209:127 (\P209:191 , \P190:127 , \G209:191 , \G190:127 , \P209:127 , \G209:127 );

  wire \G209:-1 ;

  Gij \209:-1 (\P209:127 , \G209:127 , \G126:-1 , \G209:-1 );

  Sum s210(\G209:-1 , A[210], B[210], S[210]);

  wire \P210:209 , \G210:209 ;

  PijGij \210:209 (P[210], P[209], G[210], G[209], \P210:209 , \G210:209 );

  wire \P210:207 , \G210:207 ;

  PijGij \210:207 (\P210:209 , \P208:207 , \G210:209 , \G208:207 , \P210:207 , \G210:207 );

  wire \P210:191 , \G210:191 ;

  PijGij \210:191 (\P210:207 , \P206:191 , \G210:207 , \G206:191 , \P210:191 , \G210:191 );

  wire \P210:127 , \G210:127 ;

  PijGij \210:127 (\P210:191 , \P190:127 , \G210:191 , \G190:127 , \P210:127 , \G210:127 );

  wire \G210:-1 ;

  Gij \210:-1 (\P210:127 , \G210:127 , \G126:-1 , \G210:-1 );

  Sum s211(\G210:-1 , A[211], B[211], S[211]);

  wire \P211:207 , \G211:207 ;

  PijGij \211:207 (P[211], \P210:207 , G[211], \G210:207 , \P211:207 , \G211:207 );

  wire \P211:191 , \G211:191 ;

  PijGij \211:191 (\P211:207 , \P206:191 , \G211:207 , \G206:191 , \P211:191 , \G211:191 );

  wire \P211:127 , \G211:127 ;

  PijGij \211:127 (\P211:191 , \P190:127 , \G211:191 , \G190:127 , \P211:127 , \G211:127 );

  wire \G211:-1 ;

  Gij \211:-1 (\P211:127 , \G211:127 , \G126:-1 , \G211:-1 );

  Sum s212(\G211:-1 , A[212], B[212], S[212]);

  wire \P212:211 , \G212:211 ;

  PijGij \212:211 (P[212], P[211], G[212], G[211], \P212:211 , \G212:211 );

  wire \P212:207 , \G212:207 ;

  PijGij \212:207 (\P212:211 , \P210:207 , \G212:211 , \G210:207 , \P212:207 , \G212:207 );

  wire \P212:191 , \G212:191 ;

  PijGij \212:191 (\P212:207 , \P206:191 , \G212:207 , \G206:191 , \P212:191 , \G212:191 );

  wire \P212:127 , \G212:127 ;

  PijGij \212:127 (\P212:191 , \P190:127 , \G212:191 , \G190:127 , \P212:127 , \G212:127 );

  wire \G212:-1 ;

  Gij \212:-1 (\P212:127 , \G212:127 , \G126:-1 , \G212:-1 );

  Sum s213(\G212:-1 , A[213], B[213], S[213]);

  wire \P213:211 , \G213:211 ;

  PijGij \213:211 (P[213], \P212:211 , G[213], \G212:211 , \P213:211 , \G213:211 );

  wire \P213:207 , \G213:207 ;

  PijGij \213:207 (\P213:211 , \P210:207 , \G213:211 , \G210:207 , \P213:207 , \G213:207 );

  wire \P213:191 , \G213:191 ;

  PijGij \213:191 (\P213:207 , \P206:191 , \G213:207 , \G206:191 , \P213:191 , \G213:191 );

  wire \P213:127 , \G213:127 ;

  PijGij \213:127 (\P213:191 , \P190:127 , \G213:191 , \G190:127 , \P213:127 , \G213:127 );

  wire \G213:-1 ;

  Gij \213:-1 (\P213:127 , \G213:127 , \G126:-1 , \G213:-1 );

  Sum s214(\G213:-1 , A[214], B[214], S[214]);

  wire \P214:213 , \G214:213 ;

  PijGij \214:213 (P[214], P[213], G[214], G[213], \P214:213 , \G214:213 );

  wire \P214:211 , \G214:211 ;

  PijGij \214:211 (\P214:213 , \P212:211 , \G214:213 , \G212:211 , \P214:211 , \G214:211 );

  wire \P214:207 , \G214:207 ;

  PijGij \214:207 (\P214:211 , \P210:207 , \G214:211 , \G210:207 , \P214:207 , \G214:207 );

  wire \P214:191 , \G214:191 ;

  PijGij \214:191 (\P214:207 , \P206:191 , \G214:207 , \G206:191 , \P214:191 , \G214:191 );

  wire \P214:127 , \G214:127 ;

  PijGij \214:127 (\P214:191 , \P190:127 , \G214:191 , \G190:127 , \P214:127 , \G214:127 );

  wire \G214:-1 ;

  Gij \214:-1 (\P214:127 , \G214:127 , \G126:-1 , \G214:-1 );

  Sum s215(\G214:-1 , A[215], B[215], S[215]);

  wire \P215:207 , \G215:207 ;

  PijGij \215:207 (P[215], \P214:207 , G[215], \G214:207 , \P215:207 , \G215:207 );

  wire \P215:191 , \G215:191 ;

  PijGij \215:191 (\P215:207 , \P206:191 , \G215:207 , \G206:191 , \P215:191 , \G215:191 );

  wire \P215:127 , \G215:127 ;

  PijGij \215:127 (\P215:191 , \P190:127 , \G215:191 , \G190:127 , \P215:127 , \G215:127 );

  wire \G215:-1 ;

  Gij \215:-1 (\P215:127 , \G215:127 , \G126:-1 , \G215:-1 );

  Sum s216(\G215:-1 , A[216], B[216], S[216]);

  wire \P216:215 , \G216:215 ;

  PijGij \216:215 (P[216], P[215], G[216], G[215], \P216:215 , \G216:215 );

  wire \P216:207 , \G216:207 ;

  PijGij \216:207 (\P216:215 , \P214:207 , \G216:215 , \G214:207 , \P216:207 , \G216:207 );

  wire \P216:191 , \G216:191 ;

  PijGij \216:191 (\P216:207 , \P206:191 , \G216:207 , \G206:191 , \P216:191 , \G216:191 );

  wire \P216:127 , \G216:127 ;

  PijGij \216:127 (\P216:191 , \P190:127 , \G216:191 , \G190:127 , \P216:127 , \G216:127 );

  wire \G216:-1 ;

  Gij \216:-1 (\P216:127 , \G216:127 , \G126:-1 , \G216:-1 );

  Sum s217(\G216:-1 , A[217], B[217], S[217]);

  wire \P217:215 , \G217:215 ;

  PijGij \217:215 (P[217], \P216:215 , G[217], \G216:215 , \P217:215 , \G217:215 );

  wire \P217:207 , \G217:207 ;

  PijGij \217:207 (\P217:215 , \P214:207 , \G217:215 , \G214:207 , \P217:207 , \G217:207 );

  wire \P217:191 , \G217:191 ;

  PijGij \217:191 (\P217:207 , \P206:191 , \G217:207 , \G206:191 , \P217:191 , \G217:191 );

  wire \P217:127 , \G217:127 ;

  PijGij \217:127 (\P217:191 , \P190:127 , \G217:191 , \G190:127 , \P217:127 , \G217:127 );

  wire \G217:-1 ;

  Gij \217:-1 (\P217:127 , \G217:127 , \G126:-1 , \G217:-1 );

  Sum s218(\G217:-1 , A[218], B[218], S[218]);

  wire \P218:217 , \G218:217 ;

  PijGij \218:217 (P[218], P[217], G[218], G[217], \P218:217 , \G218:217 );

  wire \P218:215 , \G218:215 ;

  PijGij \218:215 (\P218:217 , \P216:215 , \G218:217 , \G216:215 , \P218:215 , \G218:215 );

  wire \P218:207 , \G218:207 ;

  PijGij \218:207 (\P218:215 , \P214:207 , \G218:215 , \G214:207 , \P218:207 , \G218:207 );

  wire \P218:191 , \G218:191 ;

  PijGij \218:191 (\P218:207 , \P206:191 , \G218:207 , \G206:191 , \P218:191 , \G218:191 );

  wire \P218:127 , \G218:127 ;

  PijGij \218:127 (\P218:191 , \P190:127 , \G218:191 , \G190:127 , \P218:127 , \G218:127 );

  wire \G218:-1 ;

  Gij \218:-1 (\P218:127 , \G218:127 , \G126:-1 , \G218:-1 );

  Sum s219(\G218:-1 , A[219], B[219], S[219]);

  wire \P219:215 , \G219:215 ;

  PijGij \219:215 (P[219], \P218:215 , G[219], \G218:215 , \P219:215 , \G219:215 );

  wire \P219:207 , \G219:207 ;

  PijGij \219:207 (\P219:215 , \P214:207 , \G219:215 , \G214:207 , \P219:207 , \G219:207 );

  wire \P219:191 , \G219:191 ;

  PijGij \219:191 (\P219:207 , \P206:191 , \G219:207 , \G206:191 , \P219:191 , \G219:191 );

  wire \P219:127 , \G219:127 ;

  PijGij \219:127 (\P219:191 , \P190:127 , \G219:191 , \G190:127 , \P219:127 , \G219:127 );

  wire \G219:-1 ;

  Gij \219:-1 (\P219:127 , \G219:127 , \G126:-1 , \G219:-1 );

  Sum s220(\G219:-1 , A[220], B[220], S[220]);

  wire \P220:219 , \G220:219 ;

  PijGij \220:219 (P[220], P[219], G[220], G[219], \P220:219 , \G220:219 );

  wire \P220:215 , \G220:215 ;

  PijGij \220:215 (\P220:219 , \P218:215 , \G220:219 , \G218:215 , \P220:215 , \G220:215 );

  wire \P220:207 , \G220:207 ;

  PijGij \220:207 (\P220:215 , \P214:207 , \G220:215 , \G214:207 , \P220:207 , \G220:207 );

  wire \P220:191 , \G220:191 ;

  PijGij \220:191 (\P220:207 , \P206:191 , \G220:207 , \G206:191 , \P220:191 , \G220:191 );

  wire \P220:127 , \G220:127 ;

  PijGij \220:127 (\P220:191 , \P190:127 , \G220:191 , \G190:127 , \P220:127 , \G220:127 );

  wire \G220:-1 ;

  Gij \220:-1 (\P220:127 , \G220:127 , \G126:-1 , \G220:-1 );

  Sum s221(\G220:-1 , A[221], B[221], S[221]);

  wire \P221:219 , \G221:219 ;

  PijGij \221:219 (P[221], \P220:219 , G[221], \G220:219 , \P221:219 , \G221:219 );

  wire \P221:215 , \G221:215 ;

  PijGij \221:215 (\P221:219 , \P218:215 , \G221:219 , \G218:215 , \P221:215 , \G221:215 );

  wire \P221:207 , \G221:207 ;

  PijGij \221:207 (\P221:215 , \P214:207 , \G221:215 , \G214:207 , \P221:207 , \G221:207 );

  wire \P221:191 , \G221:191 ;

  PijGij \221:191 (\P221:207 , \P206:191 , \G221:207 , \G206:191 , \P221:191 , \G221:191 );

  wire \P221:127 , \G221:127 ;

  PijGij \221:127 (\P221:191 , \P190:127 , \G221:191 , \G190:127 , \P221:127 , \G221:127 );

  wire \G221:-1 ;

  Gij \221:-1 (\P221:127 , \G221:127 , \G126:-1 , \G221:-1 );

  Sum s222(\G221:-1 , A[222], B[222], S[222]);

  wire \P222:221 , \G222:221 ;

  PijGij \222:221 (P[222], P[221], G[222], G[221], \P222:221 , \G222:221 );

  wire \P222:219 , \G222:219 ;

  PijGij \222:219 (\P222:221 , \P220:219 , \G222:221 , \G220:219 , \P222:219 , \G222:219 );

  wire \P222:215 , \G222:215 ;

  PijGij \222:215 (\P222:219 , \P218:215 , \G222:219 , \G218:215 , \P222:215 , \G222:215 );

  wire \P222:207 , \G222:207 ;

  PijGij \222:207 (\P222:215 , \P214:207 , \G222:215 , \G214:207 , \P222:207 , \G222:207 );

  wire \P222:191 , \G222:191 ;

  PijGij \222:191 (\P222:207 , \P206:191 , \G222:207 , \G206:191 , \P222:191 , \G222:191 );

  wire \P222:127 , \G222:127 ;

  PijGij \222:127 (\P222:191 , \P190:127 , \G222:191 , \G190:127 , \P222:127 , \G222:127 );

  wire \G222:-1 ;

  Gij \222:-1 (\P222:127 , \G222:127 , \G126:-1 , \G222:-1 );

  Sum s223(\G222:-1 , A[223], B[223], S[223]);

  wire \P223:191 , \G223:191 ;

  PijGij \223:191 (P[223], \P222:191 , G[223], \G222:191 , \P223:191 , \G223:191 );

  wire \P223:127 , \G223:127 ;

  PijGij \223:127 (\P223:191 , \P190:127 , \G223:191 , \G190:127 , \P223:127 , \G223:127 );

  wire \G223:-1 ;

  Gij \223:-1 (\P223:127 , \G223:127 , \G126:-1 , \G223:-1 );

  Sum s224(\G223:-1 , A[224], B[224], S[224]);

  wire \P224:223 , \G224:223 ;

  PijGij \224:223 (P[224], P[223], G[224], G[223], \P224:223 , \G224:223 );

  wire \P224:191 , \G224:191 ;

  PijGij \224:191 (\P224:223 , \P222:191 , \G224:223 , \G222:191 , \P224:191 , \G224:191 );

  wire \P224:127 , \G224:127 ;

  PijGij \224:127 (\P224:191 , \P190:127 , \G224:191 , \G190:127 , \P224:127 , \G224:127 );

  wire \G224:-1 ;

  Gij \224:-1 (\P224:127 , \G224:127 , \G126:-1 , \G224:-1 );

  Sum s225(\G224:-1 , A[225], B[225], S[225]);

  wire \P225:223 , \G225:223 ;

  PijGij \225:223 (P[225], \P224:223 , G[225], \G224:223 , \P225:223 , \G225:223 );

  wire \P225:191 , \G225:191 ;

  PijGij \225:191 (\P225:223 , \P222:191 , \G225:223 , \G222:191 , \P225:191 , \G225:191 );

  wire \P225:127 , \G225:127 ;

  PijGij \225:127 (\P225:191 , \P190:127 , \G225:191 , \G190:127 , \P225:127 , \G225:127 );

  wire \G225:-1 ;

  Gij \225:-1 (\P225:127 , \G225:127 , \G126:-1 , \G225:-1 );

  Sum s226(\G225:-1 , A[226], B[226], S[226]);

  wire \P226:225 , \G226:225 ;

  PijGij \226:225 (P[226], P[225], G[226], G[225], \P226:225 , \G226:225 );

  wire \P226:223 , \G226:223 ;

  PijGij \226:223 (\P226:225 , \P224:223 , \G226:225 , \G224:223 , \P226:223 , \G226:223 );

  wire \P226:191 , \G226:191 ;

  PijGij \226:191 (\P226:223 , \P222:191 , \G226:223 , \G222:191 , \P226:191 , \G226:191 );

  wire \P226:127 , \G226:127 ;

  PijGij \226:127 (\P226:191 , \P190:127 , \G226:191 , \G190:127 , \P226:127 , \G226:127 );

  wire \G226:-1 ;

  Gij \226:-1 (\P226:127 , \G226:127 , \G126:-1 , \G226:-1 );

  Sum s227(\G226:-1 , A[227], B[227], S[227]);

  wire \P227:223 , \G227:223 ;

  PijGij \227:223 (P[227], \P226:223 , G[227], \G226:223 , \P227:223 , \G227:223 );

  wire \P227:191 , \G227:191 ;

  PijGij \227:191 (\P227:223 , \P222:191 , \G227:223 , \G222:191 , \P227:191 , \G227:191 );

  wire \P227:127 , \G227:127 ;

  PijGij \227:127 (\P227:191 , \P190:127 , \G227:191 , \G190:127 , \P227:127 , \G227:127 );

  wire \G227:-1 ;

  Gij \227:-1 (\P227:127 , \G227:127 , \G126:-1 , \G227:-1 );

  Sum s228(\G227:-1 , A[228], B[228], S[228]);

  wire \P228:227 , \G228:227 ;

  PijGij \228:227 (P[228], P[227], G[228], G[227], \P228:227 , \G228:227 );

  wire \P228:223 , \G228:223 ;

  PijGij \228:223 (\P228:227 , \P226:223 , \G228:227 , \G226:223 , \P228:223 , \G228:223 );

  wire \P228:191 , \G228:191 ;

  PijGij \228:191 (\P228:223 , \P222:191 , \G228:223 , \G222:191 , \P228:191 , \G228:191 );

  wire \P228:127 , \G228:127 ;

  PijGij \228:127 (\P228:191 , \P190:127 , \G228:191 , \G190:127 , \P228:127 , \G228:127 );

  wire \G228:-1 ;

  Gij \228:-1 (\P228:127 , \G228:127 , \G126:-1 , \G228:-1 );

  Sum s229(\G228:-1 , A[229], B[229], S[229]);

  assign Cout = (\G228:-1 & A[229]) | (\G228:-1 & B[229]) | (A[229] & B[229]);

endmodule
