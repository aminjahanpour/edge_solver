

module padder113(A, B, Cin, S, Cout);
  parameter N = 113;
  input [N-1:0] A, B;
  input Cin;
  output [N-1:0] S;
  output Cout;

  // P[i] is an alias for Pi:i, likewise G[i] is an alias for Gi:i
  wire [N-2:-1] P, G;

  assign P = {A[N-2:0] | B[N-2:0], 1'b0};
  assign G = {A[N-2:0] & B[N-2:0], Cin};

  Sum s0(G[-1], A[0], B[0], S[0]);

  wire \G0:-1 ;

  Gij \0:-1 (P[0], G[0], G[-1], \G0:-1 );

  Sum s1(\G0:-1 , A[1], B[1], S[1]);

  wire \G1:-1 ;

  Gij \1:-1 (P[1], G[1], \G0:-1 , \G1:-1 );

  Sum s2(\G1:-1 , A[2], B[2], S[2]);

  wire \P2:1 , \G2:1 ;

  PijGij \2:1 (P[2], P[1], G[2], G[1], \P2:1 , \G2:1 );

  wire \G2:-1 ;

  Gij \2:-1 (\P2:1 , \G2:1 , \G0:-1 , \G2:-1 );

  Sum s3(\G2:-1 , A[3], B[3], S[3]);

  wire \G3:-1 ;

  Gij \3:-1 (P[3], G[3], \G2:-1 , \G3:-1 );

  Sum s4(\G3:-1 , A[4], B[4], S[4]);

  wire \P4:3 , \G4:3 ;

  PijGij \4:3 (P[4], P[3], G[4], G[3], \P4:3 , \G4:3 );

  wire \G4:-1 ;

  Gij \4:-1 (\P4:3 , \G4:3 , \G2:-1 , \G4:-1 );

  Sum s5(\G4:-1 , A[5], B[5], S[5]);

  wire \P5:3 , \G5:3 ;

  PijGij \5:3 (P[5], \P4:3 , G[5], \G4:3 , \P5:3 , \G5:3 );

  wire \G5:-1 ;

  Gij \5:-1 (\P5:3 , \G5:3 , \G2:-1 , \G5:-1 );

  Sum s6(\G5:-1 , A[6], B[6], S[6]);

  wire \P6:5 , \G6:5 ;

  PijGij \6:5 (P[6], P[5], G[6], G[5], \P6:5 , \G6:5 );

  wire \P6:3 , \G6:3 ;

  PijGij \6:3 (\P6:5 , \P4:3 , \G6:5 , \G4:3 , \P6:3 , \G6:3 );

  wire \G6:-1 ;

  Gij \6:-1 (\P6:3 , \G6:3 , \G2:-1 , \G6:-1 );

  Sum s7(\G6:-1 , A[7], B[7], S[7]);

  wire \G7:-1 ;

  Gij \7:-1 (P[7], G[7], \G6:-1 , \G7:-1 );

  Sum s8(\G7:-1 , A[8], B[8], S[8]);

  wire \P8:7 , \G8:7 ;

  PijGij \8:7 (P[8], P[7], G[8], G[7], \P8:7 , \G8:7 );

  wire \G8:-1 ;

  Gij \8:-1 (\P8:7 , \G8:7 , \G6:-1 , \G8:-1 );

  Sum s9(\G8:-1 , A[9], B[9], S[9]);

  wire \P9:7 , \G9:7 ;

  PijGij \9:7 (P[9], \P8:7 , G[9], \G8:7 , \P9:7 , \G9:7 );

  wire \G9:-1 ;

  Gij \9:-1 (\P9:7 , \G9:7 , \G6:-1 , \G9:-1 );

  Sum s10(\G9:-1 , A[10], B[10], S[10]);

  wire \P10:9 , \G10:9 ;

  PijGij \10:9 (P[10], P[9], G[10], G[9], \P10:9 , \G10:9 );

  wire \P10:7 , \G10:7 ;

  PijGij \10:7 (\P10:9 , \P8:7 , \G10:9 , \G8:7 , \P10:7 , \G10:7 );

  wire \G10:-1 ;

  Gij \10:-1 (\P10:7 , \G10:7 , \G6:-1 , \G10:-1 );

  Sum s11(\G10:-1 , A[11], B[11], S[11]);

  wire \P11:7 , \G11:7 ;

  PijGij \11:7 (P[11], \P10:7 , G[11], \G10:7 , \P11:7 , \G11:7 );

  wire \G11:-1 ;

  Gij \11:-1 (\P11:7 , \G11:7 , \G6:-1 , \G11:-1 );

  Sum s12(\G11:-1 , A[12], B[12], S[12]);

  wire \P12:11 , \G12:11 ;

  PijGij \12:11 (P[12], P[11], G[12], G[11], \P12:11 , \G12:11 );

  wire \P12:7 , \G12:7 ;

  PijGij \12:7 (\P12:11 , \P10:7 , \G12:11 , \G10:7 , \P12:7 , \G12:7 );

  wire \G12:-1 ;

  Gij \12:-1 (\P12:7 , \G12:7 , \G6:-1 , \G12:-1 );

  Sum s13(\G12:-1 , A[13], B[13], S[13]);

  wire \P13:11 , \G13:11 ;

  PijGij \13:11 (P[13], \P12:11 , G[13], \G12:11 , \P13:11 , \G13:11 );

  wire \P13:7 , \G13:7 ;

  PijGij \13:7 (\P13:11 , \P10:7 , \G13:11 , \G10:7 , \P13:7 , \G13:7 );

  wire \G13:-1 ;

  Gij \13:-1 (\P13:7 , \G13:7 , \G6:-1 , \G13:-1 );

  Sum s14(\G13:-1 , A[14], B[14], S[14]);

  wire \P14:13 , \G14:13 ;

  PijGij \14:13 (P[14], P[13], G[14], G[13], \P14:13 , \G14:13 );

  wire \P14:11 , \G14:11 ;

  PijGij \14:11 (\P14:13 , \P12:11 , \G14:13 , \G12:11 , \P14:11 , \G14:11 );

  wire \P14:7 , \G14:7 ;

  PijGij \14:7 (\P14:11 , \P10:7 , \G14:11 , \G10:7 , \P14:7 , \G14:7 );

  wire \G14:-1 ;

  Gij \14:-1 (\P14:7 , \G14:7 , \G6:-1 , \G14:-1 );

  Sum s15(\G14:-1 , A[15], B[15], S[15]);

  wire \G15:-1 ;

  Gij \15:-1 (P[15], G[15], \G14:-1 , \G15:-1 );

  Sum s16(\G15:-1 , A[16], B[16], S[16]);

  wire \P16:15 , \G16:15 ;

  PijGij \16:15 (P[16], P[15], G[16], G[15], \P16:15 , \G16:15 );

  wire \G16:-1 ;

  Gij \16:-1 (\P16:15 , \G16:15 , \G14:-1 , \G16:-1 );

  Sum s17(\G16:-1 , A[17], B[17], S[17]);

  wire \P17:15 , \G17:15 ;

  PijGij \17:15 (P[17], \P16:15 , G[17], \G16:15 , \P17:15 , \G17:15 );

  wire \G17:-1 ;

  Gij \17:-1 (\P17:15 , \G17:15 , \G14:-1 , \G17:-1 );

  Sum s18(\G17:-1 , A[18], B[18], S[18]);

  wire \P18:17 , \G18:17 ;

  PijGij \18:17 (P[18], P[17], G[18], G[17], \P18:17 , \G18:17 );

  wire \P18:15 , \G18:15 ;

  PijGij \18:15 (\P18:17 , \P16:15 , \G18:17 , \G16:15 , \P18:15 , \G18:15 );

  wire \G18:-1 ;

  Gij \18:-1 (\P18:15 , \G18:15 , \G14:-1 , \G18:-1 );

  Sum s19(\G18:-1 , A[19], B[19], S[19]);

  wire \P19:15 , \G19:15 ;

  PijGij \19:15 (P[19], \P18:15 , G[19], \G18:15 , \P19:15 , \G19:15 );

  wire \G19:-1 ;

  Gij \19:-1 (\P19:15 , \G19:15 , \G14:-1 , \G19:-1 );

  Sum s20(\G19:-1 , A[20], B[20], S[20]);

  wire \P20:19 , \G20:19 ;

  PijGij \20:19 (P[20], P[19], G[20], G[19], \P20:19 , \G20:19 );

  wire \P20:15 , \G20:15 ;

  PijGij \20:15 (\P20:19 , \P18:15 , \G20:19 , \G18:15 , \P20:15 , \G20:15 );

  wire \G20:-1 ;

  Gij \20:-1 (\P20:15 , \G20:15 , \G14:-1 , \G20:-1 );

  Sum s21(\G20:-1 , A[21], B[21], S[21]);

  wire \P21:19 , \G21:19 ;

  PijGij \21:19 (P[21], \P20:19 , G[21], \G20:19 , \P21:19 , \G21:19 );

  wire \P21:15 , \G21:15 ;

  PijGij \21:15 (\P21:19 , \P18:15 , \G21:19 , \G18:15 , \P21:15 , \G21:15 );

  wire \G21:-1 ;

  Gij \21:-1 (\P21:15 , \G21:15 , \G14:-1 , \G21:-1 );

  Sum s22(\G21:-1 , A[22], B[22], S[22]);

  wire \P22:21 , \G22:21 ;

  PijGij \22:21 (P[22], P[21], G[22], G[21], \P22:21 , \G22:21 );

  wire \P22:19 , \G22:19 ;

  PijGij \22:19 (\P22:21 , \P20:19 , \G22:21 , \G20:19 , \P22:19 , \G22:19 );

  wire \P22:15 , \G22:15 ;

  PijGij \22:15 (\P22:19 , \P18:15 , \G22:19 , \G18:15 , \P22:15 , \G22:15 );

  wire \G22:-1 ;

  Gij \22:-1 (\P22:15 , \G22:15 , \G14:-1 , \G22:-1 );

  Sum s23(\G22:-1 , A[23], B[23], S[23]);

  wire \P23:15 , \G23:15 ;

  PijGij \23:15 (P[23], \P22:15 , G[23], \G22:15 , \P23:15 , \G23:15 );

  wire \G23:-1 ;

  Gij \23:-1 (\P23:15 , \G23:15 , \G14:-1 , \G23:-1 );

  Sum s24(\G23:-1 , A[24], B[24], S[24]);

  wire \P24:23 , \G24:23 ;

  PijGij \24:23 (P[24], P[23], G[24], G[23], \P24:23 , \G24:23 );

  wire \P24:15 , \G24:15 ;

  PijGij \24:15 (\P24:23 , \P22:15 , \G24:23 , \G22:15 , \P24:15 , \G24:15 );

  wire \G24:-1 ;

  Gij \24:-1 (\P24:15 , \G24:15 , \G14:-1 , \G24:-1 );

  Sum s25(\G24:-1 , A[25], B[25], S[25]);

  wire \P25:23 , \G25:23 ;

  PijGij \25:23 (P[25], \P24:23 , G[25], \G24:23 , \P25:23 , \G25:23 );

  wire \P25:15 , \G25:15 ;

  PijGij \25:15 (\P25:23 , \P22:15 , \G25:23 , \G22:15 , \P25:15 , \G25:15 );

  wire \G25:-1 ;

  Gij \25:-1 (\P25:15 , \G25:15 , \G14:-1 , \G25:-1 );

  Sum s26(\G25:-1 , A[26], B[26], S[26]);

  wire \P26:25 , \G26:25 ;

  PijGij \26:25 (P[26], P[25], G[26], G[25], \P26:25 , \G26:25 );

  wire \P26:23 , \G26:23 ;

  PijGij \26:23 (\P26:25 , \P24:23 , \G26:25 , \G24:23 , \P26:23 , \G26:23 );

  wire \P26:15 , \G26:15 ;

  PijGij \26:15 (\P26:23 , \P22:15 , \G26:23 , \G22:15 , \P26:15 , \G26:15 );

  wire \G26:-1 ;

  Gij \26:-1 (\P26:15 , \G26:15 , \G14:-1 , \G26:-1 );

  Sum s27(\G26:-1 , A[27], B[27], S[27]);

  wire \P27:23 , \G27:23 ;

  PijGij \27:23 (P[27], \P26:23 , G[27], \G26:23 , \P27:23 , \G27:23 );

  wire \P27:15 , \G27:15 ;

  PijGij \27:15 (\P27:23 , \P22:15 , \G27:23 , \G22:15 , \P27:15 , \G27:15 );

  wire \G27:-1 ;

  Gij \27:-1 (\P27:15 , \G27:15 , \G14:-1 , \G27:-1 );

  Sum s28(\G27:-1 , A[28], B[28], S[28]);

  wire \P28:27 , \G28:27 ;

  PijGij \28:27 (P[28], P[27], G[28], G[27], \P28:27 , \G28:27 );

  wire \P28:23 , \G28:23 ;

  PijGij \28:23 (\P28:27 , \P26:23 , \G28:27 , \G26:23 , \P28:23 , \G28:23 );

  wire \P28:15 , \G28:15 ;

  PijGij \28:15 (\P28:23 , \P22:15 , \G28:23 , \G22:15 , \P28:15 , \G28:15 );

  wire \G28:-1 ;

  Gij \28:-1 (\P28:15 , \G28:15 , \G14:-1 , \G28:-1 );

  Sum s29(\G28:-1 , A[29], B[29], S[29]);

  wire \P29:27 , \G29:27 ;

  PijGij \29:27 (P[29], \P28:27 , G[29], \G28:27 , \P29:27 , \G29:27 );

  wire \P29:23 , \G29:23 ;

  PijGij \29:23 (\P29:27 , \P26:23 , \G29:27 , \G26:23 , \P29:23 , \G29:23 );

  wire \P29:15 , \G29:15 ;

  PijGij \29:15 (\P29:23 , \P22:15 , \G29:23 , \G22:15 , \P29:15 , \G29:15 );

  wire \G29:-1 ;

  Gij \29:-1 (\P29:15 , \G29:15 , \G14:-1 , \G29:-1 );

  Sum s30(\G29:-1 , A[30], B[30], S[30]);

  wire \P30:29 , \G30:29 ;

  PijGij \30:29 (P[30], P[29], G[30], G[29], \P30:29 , \G30:29 );

  wire \P30:27 , \G30:27 ;

  PijGij \30:27 (\P30:29 , \P28:27 , \G30:29 , \G28:27 , \P30:27 , \G30:27 );

  wire \P30:23 , \G30:23 ;

  PijGij \30:23 (\P30:27 , \P26:23 , \G30:27 , \G26:23 , \P30:23 , \G30:23 );

  wire \P30:15 , \G30:15 ;

  PijGij \30:15 (\P30:23 , \P22:15 , \G30:23 , \G22:15 , \P30:15 , \G30:15 );

  wire \G30:-1 ;

  Gij \30:-1 (\P30:15 , \G30:15 , \G14:-1 , \G30:-1 );

  Sum s31(\G30:-1 , A[31], B[31], S[31]);

  wire \G31:-1 ;

  Gij \31:-1 (P[31], G[31], \G30:-1 , \G31:-1 );

  Sum s32(\G31:-1 , A[32], B[32], S[32]);

  wire \P32:31 , \G32:31 ;

  PijGij \32:31 (P[32], P[31], G[32], G[31], \P32:31 , \G32:31 );

  wire \G32:-1 ;

  Gij \32:-1 (\P32:31 , \G32:31 , \G30:-1 , \G32:-1 );

  Sum s33(\G32:-1 , A[33], B[33], S[33]);

  wire \P33:31 , \G33:31 ;

  PijGij \33:31 (P[33], \P32:31 , G[33], \G32:31 , \P33:31 , \G33:31 );

  wire \G33:-1 ;

  Gij \33:-1 (\P33:31 , \G33:31 , \G30:-1 , \G33:-1 );

  Sum s34(\G33:-1 , A[34], B[34], S[34]);

  wire \P34:33 , \G34:33 ;

  PijGij \34:33 (P[34], P[33], G[34], G[33], \P34:33 , \G34:33 );

  wire \P34:31 , \G34:31 ;

  PijGij \34:31 (\P34:33 , \P32:31 , \G34:33 , \G32:31 , \P34:31 , \G34:31 );

  wire \G34:-1 ;

  Gij \34:-1 (\P34:31 , \G34:31 , \G30:-1 , \G34:-1 );

  Sum s35(\G34:-1 , A[35], B[35], S[35]);

  wire \P35:31 , \G35:31 ;

  PijGij \35:31 (P[35], \P34:31 , G[35], \G34:31 , \P35:31 , \G35:31 );

  wire \G35:-1 ;

  Gij \35:-1 (\P35:31 , \G35:31 , \G30:-1 , \G35:-1 );

  Sum s36(\G35:-1 , A[36], B[36], S[36]);

  wire \P36:35 , \G36:35 ;

  PijGij \36:35 (P[36], P[35], G[36], G[35], \P36:35 , \G36:35 );

  wire \P36:31 , \G36:31 ;

  PijGij \36:31 (\P36:35 , \P34:31 , \G36:35 , \G34:31 , \P36:31 , \G36:31 );

  wire \G36:-1 ;

  Gij \36:-1 (\P36:31 , \G36:31 , \G30:-1 , \G36:-1 );

  Sum s37(\G36:-1 , A[37], B[37], S[37]);

  wire \P37:35 , \G37:35 ;

  PijGij \37:35 (P[37], \P36:35 , G[37], \G36:35 , \P37:35 , \G37:35 );

  wire \P37:31 , \G37:31 ;

  PijGij \37:31 (\P37:35 , \P34:31 , \G37:35 , \G34:31 , \P37:31 , \G37:31 );

  wire \G37:-1 ;

  Gij \37:-1 (\P37:31 , \G37:31 , \G30:-1 , \G37:-1 );

  Sum s38(\G37:-1 , A[38], B[38], S[38]);

  wire \P38:37 , \G38:37 ;

  PijGij \38:37 (P[38], P[37], G[38], G[37], \P38:37 , \G38:37 );

  wire \P38:35 , \G38:35 ;

  PijGij \38:35 (\P38:37 , \P36:35 , \G38:37 , \G36:35 , \P38:35 , \G38:35 );

  wire \P38:31 , \G38:31 ;

  PijGij \38:31 (\P38:35 , \P34:31 , \G38:35 , \G34:31 , \P38:31 , \G38:31 );

  wire \G38:-1 ;

  Gij \38:-1 (\P38:31 , \G38:31 , \G30:-1 , \G38:-1 );

  Sum s39(\G38:-1 , A[39], B[39], S[39]);

  wire \P39:31 , \G39:31 ;

  PijGij \39:31 (P[39], \P38:31 , G[39], \G38:31 , \P39:31 , \G39:31 );

  wire \G39:-1 ;

  Gij \39:-1 (\P39:31 , \G39:31 , \G30:-1 , \G39:-1 );

  Sum s40(\G39:-1 , A[40], B[40], S[40]);

  wire \P40:39 , \G40:39 ;

  PijGij \40:39 (P[40], P[39], G[40], G[39], \P40:39 , \G40:39 );

  wire \P40:31 , \G40:31 ;

  PijGij \40:31 (\P40:39 , \P38:31 , \G40:39 , \G38:31 , \P40:31 , \G40:31 );

  wire \G40:-1 ;

  Gij \40:-1 (\P40:31 , \G40:31 , \G30:-1 , \G40:-1 );

  Sum s41(\G40:-1 , A[41], B[41], S[41]);

  wire \P41:39 , \G41:39 ;

  PijGij \41:39 (P[41], \P40:39 , G[41], \G40:39 , \P41:39 , \G41:39 );

  wire \P41:31 , \G41:31 ;

  PijGij \41:31 (\P41:39 , \P38:31 , \G41:39 , \G38:31 , \P41:31 , \G41:31 );

  wire \G41:-1 ;

  Gij \41:-1 (\P41:31 , \G41:31 , \G30:-1 , \G41:-1 );

  Sum s42(\G41:-1 , A[42], B[42], S[42]);

  wire \P42:41 , \G42:41 ;

  PijGij \42:41 (P[42], P[41], G[42], G[41], \P42:41 , \G42:41 );

  wire \P42:39 , \G42:39 ;

  PijGij \42:39 (\P42:41 , \P40:39 , \G42:41 , \G40:39 , \P42:39 , \G42:39 );

  wire \P42:31 , \G42:31 ;

  PijGij \42:31 (\P42:39 , \P38:31 , \G42:39 , \G38:31 , \P42:31 , \G42:31 );

  wire \G42:-1 ;

  Gij \42:-1 (\P42:31 , \G42:31 , \G30:-1 , \G42:-1 );

  Sum s43(\G42:-1 , A[43], B[43], S[43]);

  wire \P43:39 , \G43:39 ;

  PijGij \43:39 (P[43], \P42:39 , G[43], \G42:39 , \P43:39 , \G43:39 );

  wire \P43:31 , \G43:31 ;

  PijGij \43:31 (\P43:39 , \P38:31 , \G43:39 , \G38:31 , \P43:31 , \G43:31 );

  wire \G43:-1 ;

  Gij \43:-1 (\P43:31 , \G43:31 , \G30:-1 , \G43:-1 );

  Sum s44(\G43:-1 , A[44], B[44], S[44]);

  wire \P44:43 , \G44:43 ;

  PijGij \44:43 (P[44], P[43], G[44], G[43], \P44:43 , \G44:43 );

  wire \P44:39 , \G44:39 ;

  PijGij \44:39 (\P44:43 , \P42:39 , \G44:43 , \G42:39 , \P44:39 , \G44:39 );

  wire \P44:31 , \G44:31 ;

  PijGij \44:31 (\P44:39 , \P38:31 , \G44:39 , \G38:31 , \P44:31 , \G44:31 );

  wire \G44:-1 ;

  Gij \44:-1 (\P44:31 , \G44:31 , \G30:-1 , \G44:-1 );

  Sum s45(\G44:-1 , A[45], B[45], S[45]);

  wire \P45:43 , \G45:43 ;

  PijGij \45:43 (P[45], \P44:43 , G[45], \G44:43 , \P45:43 , \G45:43 );

  wire \P45:39 , \G45:39 ;

  PijGij \45:39 (\P45:43 , \P42:39 , \G45:43 , \G42:39 , \P45:39 , \G45:39 );

  wire \P45:31 , \G45:31 ;

  PijGij \45:31 (\P45:39 , \P38:31 , \G45:39 , \G38:31 , \P45:31 , \G45:31 );

  wire \G45:-1 ;

  Gij \45:-1 (\P45:31 , \G45:31 , \G30:-1 , \G45:-1 );

  Sum s46(\G45:-1 , A[46], B[46], S[46]);

  wire \P46:45 , \G46:45 ;

  PijGij \46:45 (P[46], P[45], G[46], G[45], \P46:45 , \G46:45 );

  wire \P46:43 , \G46:43 ;

  PijGij \46:43 (\P46:45 , \P44:43 , \G46:45 , \G44:43 , \P46:43 , \G46:43 );

  wire \P46:39 , \G46:39 ;

  PijGij \46:39 (\P46:43 , \P42:39 , \G46:43 , \G42:39 , \P46:39 , \G46:39 );

  wire \P46:31 , \G46:31 ;

  PijGij \46:31 (\P46:39 , \P38:31 , \G46:39 , \G38:31 , \P46:31 , \G46:31 );

  wire \G46:-1 ;

  Gij \46:-1 (\P46:31 , \G46:31 , \G30:-1 , \G46:-1 );

  Sum s47(\G46:-1 , A[47], B[47], S[47]);

  wire \P47:31 , \G47:31 ;

  PijGij \47:31 (P[47], \P46:31 , G[47], \G46:31 , \P47:31 , \G47:31 );

  wire \G47:-1 ;

  Gij \47:-1 (\P47:31 , \G47:31 , \G30:-1 , \G47:-1 );

  Sum s48(\G47:-1 , A[48], B[48], S[48]);

  wire \P48:47 , \G48:47 ;

  PijGij \48:47 (P[48], P[47], G[48], G[47], \P48:47 , \G48:47 );

  wire \P48:31 , \G48:31 ;

  PijGij \48:31 (\P48:47 , \P46:31 , \G48:47 , \G46:31 , \P48:31 , \G48:31 );

  wire \G48:-1 ;

  Gij \48:-1 (\P48:31 , \G48:31 , \G30:-1 , \G48:-1 );

  Sum s49(\G48:-1 , A[49], B[49], S[49]);

  wire \P49:47 , \G49:47 ;

  PijGij \49:47 (P[49], \P48:47 , G[49], \G48:47 , \P49:47 , \G49:47 );

  wire \P49:31 , \G49:31 ;

  PijGij \49:31 (\P49:47 , \P46:31 , \G49:47 , \G46:31 , \P49:31 , \G49:31 );

  wire \G49:-1 ;

  Gij \49:-1 (\P49:31 , \G49:31 , \G30:-1 , \G49:-1 );

  Sum s50(\G49:-1 , A[50], B[50], S[50]);

  wire \P50:49 , \G50:49 ;

  PijGij \50:49 (P[50], P[49], G[50], G[49], \P50:49 , \G50:49 );

  wire \P50:47 , \G50:47 ;

  PijGij \50:47 (\P50:49 , \P48:47 , \G50:49 , \G48:47 , \P50:47 , \G50:47 );

  wire \P50:31 , \G50:31 ;

  PijGij \50:31 (\P50:47 , \P46:31 , \G50:47 , \G46:31 , \P50:31 , \G50:31 );

  wire \G50:-1 ;

  Gij \50:-1 (\P50:31 , \G50:31 , \G30:-1 , \G50:-1 );

  Sum s51(\G50:-1 , A[51], B[51], S[51]);

  wire \P51:47 , \G51:47 ;

  PijGij \51:47 (P[51], \P50:47 , G[51], \G50:47 , \P51:47 , \G51:47 );

  wire \P51:31 , \G51:31 ;

  PijGij \51:31 (\P51:47 , \P46:31 , \G51:47 , \G46:31 , \P51:31 , \G51:31 );

  wire \G51:-1 ;

  Gij \51:-1 (\P51:31 , \G51:31 , \G30:-1 , \G51:-1 );

  Sum s52(\G51:-1 , A[52], B[52], S[52]);

  wire \P52:51 , \G52:51 ;

  PijGij \52:51 (P[52], P[51], G[52], G[51], \P52:51 , \G52:51 );

  wire \P52:47 , \G52:47 ;

  PijGij \52:47 (\P52:51 , \P50:47 , \G52:51 , \G50:47 , \P52:47 , \G52:47 );

  wire \P52:31 , \G52:31 ;

  PijGij \52:31 (\P52:47 , \P46:31 , \G52:47 , \G46:31 , \P52:31 , \G52:31 );

  wire \G52:-1 ;

  Gij \52:-1 (\P52:31 , \G52:31 , \G30:-1 , \G52:-1 );

  Sum s53(\G52:-1 , A[53], B[53], S[53]);

  wire \P53:51 , \G53:51 ;

  PijGij \53:51 (P[53], \P52:51 , G[53], \G52:51 , \P53:51 , \G53:51 );

  wire \P53:47 , \G53:47 ;

  PijGij \53:47 (\P53:51 , \P50:47 , \G53:51 , \G50:47 , \P53:47 , \G53:47 );

  wire \P53:31 , \G53:31 ;

  PijGij \53:31 (\P53:47 , \P46:31 , \G53:47 , \G46:31 , \P53:31 , \G53:31 );

  wire \G53:-1 ;

  Gij \53:-1 (\P53:31 , \G53:31 , \G30:-1 , \G53:-1 );

  Sum s54(\G53:-1 , A[54], B[54], S[54]);

  wire \P54:53 , \G54:53 ;

  PijGij \54:53 (P[54], P[53], G[54], G[53], \P54:53 , \G54:53 );

  wire \P54:51 , \G54:51 ;

  PijGij \54:51 (\P54:53 , \P52:51 , \G54:53 , \G52:51 , \P54:51 , \G54:51 );

  wire \P54:47 , \G54:47 ;

  PijGij \54:47 (\P54:51 , \P50:47 , \G54:51 , \G50:47 , \P54:47 , \G54:47 );

  wire \P54:31 , \G54:31 ;

  PijGij \54:31 (\P54:47 , \P46:31 , \G54:47 , \G46:31 , \P54:31 , \G54:31 );

  wire \G54:-1 ;

  Gij \54:-1 (\P54:31 , \G54:31 , \G30:-1 , \G54:-1 );

  Sum s55(\G54:-1 , A[55], B[55], S[55]);

  wire \P55:47 , \G55:47 ;

  PijGij \55:47 (P[55], \P54:47 , G[55], \G54:47 , \P55:47 , \G55:47 );

  wire \P55:31 , \G55:31 ;

  PijGij \55:31 (\P55:47 , \P46:31 , \G55:47 , \G46:31 , \P55:31 , \G55:31 );

  wire \G55:-1 ;

  Gij \55:-1 (\P55:31 , \G55:31 , \G30:-1 , \G55:-1 );

  Sum s56(\G55:-1 , A[56], B[56], S[56]);

  wire \P56:55 , \G56:55 ;

  PijGij \56:55 (P[56], P[55], G[56], G[55], \P56:55 , \G56:55 );

  wire \P56:47 , \G56:47 ;

  PijGij \56:47 (\P56:55 , \P54:47 , \G56:55 , \G54:47 , \P56:47 , \G56:47 );

  wire \P56:31 , \G56:31 ;

  PijGij \56:31 (\P56:47 , \P46:31 , \G56:47 , \G46:31 , \P56:31 , \G56:31 );

  wire \G56:-1 ;

  Gij \56:-1 (\P56:31 , \G56:31 , \G30:-1 , \G56:-1 );

  Sum s57(\G56:-1 , A[57], B[57], S[57]);

  wire \P57:55 , \G57:55 ;

  PijGij \57:55 (P[57], \P56:55 , G[57], \G56:55 , \P57:55 , \G57:55 );

  wire \P57:47 , \G57:47 ;

  PijGij \57:47 (\P57:55 , \P54:47 , \G57:55 , \G54:47 , \P57:47 , \G57:47 );

  wire \P57:31 , \G57:31 ;

  PijGij \57:31 (\P57:47 , \P46:31 , \G57:47 , \G46:31 , \P57:31 , \G57:31 );

  wire \G57:-1 ;

  Gij \57:-1 (\P57:31 , \G57:31 , \G30:-1 , \G57:-1 );

  Sum s58(\G57:-1 , A[58], B[58], S[58]);

  wire \P58:57 , \G58:57 ;

  PijGij \58:57 (P[58], P[57], G[58], G[57], \P58:57 , \G58:57 );

  wire \P58:55 , \G58:55 ;

  PijGij \58:55 (\P58:57 , \P56:55 , \G58:57 , \G56:55 , \P58:55 , \G58:55 );

  wire \P58:47 , \G58:47 ;

  PijGij \58:47 (\P58:55 , \P54:47 , \G58:55 , \G54:47 , \P58:47 , \G58:47 );

  wire \P58:31 , \G58:31 ;

  PijGij \58:31 (\P58:47 , \P46:31 , \G58:47 , \G46:31 , \P58:31 , \G58:31 );

  wire \G58:-1 ;

  Gij \58:-1 (\P58:31 , \G58:31 , \G30:-1 , \G58:-1 );

  Sum s59(\G58:-1 , A[59], B[59], S[59]);

  wire \P59:55 , \G59:55 ;

  PijGij \59:55 (P[59], \P58:55 , G[59], \G58:55 , \P59:55 , \G59:55 );

  wire \P59:47 , \G59:47 ;

  PijGij \59:47 (\P59:55 , \P54:47 , \G59:55 , \G54:47 , \P59:47 , \G59:47 );

  wire \P59:31 , \G59:31 ;

  PijGij \59:31 (\P59:47 , \P46:31 , \G59:47 , \G46:31 , \P59:31 , \G59:31 );

  wire \G59:-1 ;

  Gij \59:-1 (\P59:31 , \G59:31 , \G30:-1 , \G59:-1 );

  Sum s60(\G59:-1 , A[60], B[60], S[60]);

  wire \P60:59 , \G60:59 ;

  PijGij \60:59 (P[60], P[59], G[60], G[59], \P60:59 , \G60:59 );

  wire \P60:55 , \G60:55 ;

  PijGij \60:55 (\P60:59 , \P58:55 , \G60:59 , \G58:55 , \P60:55 , \G60:55 );

  wire \P60:47 , \G60:47 ;

  PijGij \60:47 (\P60:55 , \P54:47 , \G60:55 , \G54:47 , \P60:47 , \G60:47 );

  wire \P60:31 , \G60:31 ;

  PijGij \60:31 (\P60:47 , \P46:31 , \G60:47 , \G46:31 , \P60:31 , \G60:31 );

  wire \G60:-1 ;

  Gij \60:-1 (\P60:31 , \G60:31 , \G30:-1 , \G60:-1 );

  Sum s61(\G60:-1 , A[61], B[61], S[61]);

  wire \P61:59 , \G61:59 ;

  PijGij \61:59 (P[61], \P60:59 , G[61], \G60:59 , \P61:59 , \G61:59 );

  wire \P61:55 , \G61:55 ;

  PijGij \61:55 (\P61:59 , \P58:55 , \G61:59 , \G58:55 , \P61:55 , \G61:55 );

  wire \P61:47 , \G61:47 ;

  PijGij \61:47 (\P61:55 , \P54:47 , \G61:55 , \G54:47 , \P61:47 , \G61:47 );

  wire \P61:31 , \G61:31 ;

  PijGij \61:31 (\P61:47 , \P46:31 , \G61:47 , \G46:31 , \P61:31 , \G61:31 );

  wire \G61:-1 ;

  Gij \61:-1 (\P61:31 , \G61:31 , \G30:-1 , \G61:-1 );

  Sum s62(\G61:-1 , A[62], B[62], S[62]);

  wire \P62:61 , \G62:61 ;

  PijGij \62:61 (P[62], P[61], G[62], G[61], \P62:61 , \G62:61 );

  wire \P62:59 , \G62:59 ;

  PijGij \62:59 (\P62:61 , \P60:59 , \G62:61 , \G60:59 , \P62:59 , \G62:59 );

  wire \P62:55 , \G62:55 ;

  PijGij \62:55 (\P62:59 , \P58:55 , \G62:59 , \G58:55 , \P62:55 , \G62:55 );

  wire \P62:47 , \G62:47 ;

  PijGij \62:47 (\P62:55 , \P54:47 , \G62:55 , \G54:47 , \P62:47 , \G62:47 );

  wire \P62:31 , \G62:31 ;

  PijGij \62:31 (\P62:47 , \P46:31 , \G62:47 , \G46:31 , \P62:31 , \G62:31 );

  wire \G62:-1 ;

  Gij \62:-1 (\P62:31 , \G62:31 , \G30:-1 , \G62:-1 );

  Sum s63(\G62:-1 , A[63], B[63], S[63]);

  wire \G63:-1 ;

  Gij \63:-1 (P[63], G[63], \G62:-1 , \G63:-1 );

  Sum s64(\G63:-1 , A[64], B[64], S[64]);

  wire \P64:63 , \G64:63 ;

  PijGij \64:63 (P[64], P[63], G[64], G[63], \P64:63 , \G64:63 );

  wire \G64:-1 ;

  Gij \64:-1 (\P64:63 , \G64:63 , \G62:-1 , \G64:-1 );

  Sum s65(\G64:-1 , A[65], B[65], S[65]);

  wire \P65:63 , \G65:63 ;

  PijGij \65:63 (P[65], \P64:63 , G[65], \G64:63 , \P65:63 , \G65:63 );

  wire \G65:-1 ;

  Gij \65:-1 (\P65:63 , \G65:63 , \G62:-1 , \G65:-1 );

  Sum s66(\G65:-1 , A[66], B[66], S[66]);

  wire \P66:65 , \G66:65 ;

  PijGij \66:65 (P[66], P[65], G[66], G[65], \P66:65 , \G66:65 );

  wire \P66:63 , \G66:63 ;

  PijGij \66:63 (\P66:65 , \P64:63 , \G66:65 , \G64:63 , \P66:63 , \G66:63 );

  wire \G66:-1 ;

  Gij \66:-1 (\P66:63 , \G66:63 , \G62:-1 , \G66:-1 );

  Sum s67(\G66:-1 , A[67], B[67], S[67]);

  wire \P67:63 , \G67:63 ;

  PijGij \67:63 (P[67], \P66:63 , G[67], \G66:63 , \P67:63 , \G67:63 );

  wire \G67:-1 ;

  Gij \67:-1 (\P67:63 , \G67:63 , \G62:-1 , \G67:-1 );

  Sum s68(\G67:-1 , A[68], B[68], S[68]);

  wire \P68:67 , \G68:67 ;

  PijGij \68:67 (P[68], P[67], G[68], G[67], \P68:67 , \G68:67 );

  wire \P68:63 , \G68:63 ;

  PijGij \68:63 (\P68:67 , \P66:63 , \G68:67 , \G66:63 , \P68:63 , \G68:63 );

  wire \G68:-1 ;

  Gij \68:-1 (\P68:63 , \G68:63 , \G62:-1 , \G68:-1 );

  Sum s69(\G68:-1 , A[69], B[69], S[69]);

  wire \P69:67 , \G69:67 ;

  PijGij \69:67 (P[69], \P68:67 , G[69], \G68:67 , \P69:67 , \G69:67 );

  wire \P69:63 , \G69:63 ;

  PijGij \69:63 (\P69:67 , \P66:63 , \G69:67 , \G66:63 , \P69:63 , \G69:63 );

  wire \G69:-1 ;

  Gij \69:-1 (\P69:63 , \G69:63 , \G62:-1 , \G69:-1 );

  Sum s70(\G69:-1 , A[70], B[70], S[70]);

  wire \P70:69 , \G70:69 ;

  PijGij \70:69 (P[70], P[69], G[70], G[69], \P70:69 , \G70:69 );

  wire \P70:67 , \G70:67 ;

  PijGij \70:67 (\P70:69 , \P68:67 , \G70:69 , \G68:67 , \P70:67 , \G70:67 );

  wire \P70:63 , \G70:63 ;

  PijGij \70:63 (\P70:67 , \P66:63 , \G70:67 , \G66:63 , \P70:63 , \G70:63 );

  wire \G70:-1 ;

  Gij \70:-1 (\P70:63 , \G70:63 , \G62:-1 , \G70:-1 );

  Sum s71(\G70:-1 , A[71], B[71], S[71]);

  wire \P71:63 , \G71:63 ;

  PijGij \71:63 (P[71], \P70:63 , G[71], \G70:63 , \P71:63 , \G71:63 );

  wire \G71:-1 ;

  Gij \71:-1 (\P71:63 , \G71:63 , \G62:-1 , \G71:-1 );

  Sum s72(\G71:-1 , A[72], B[72], S[72]);

  wire \P72:71 , \G72:71 ;

  PijGij \72:71 (P[72], P[71], G[72], G[71], \P72:71 , \G72:71 );

  wire \P72:63 , \G72:63 ;

  PijGij \72:63 (\P72:71 , \P70:63 , \G72:71 , \G70:63 , \P72:63 , \G72:63 );

  wire \G72:-1 ;

  Gij \72:-1 (\P72:63 , \G72:63 , \G62:-1 , \G72:-1 );

  Sum s73(\G72:-1 , A[73], B[73], S[73]);

  wire \P73:71 , \G73:71 ;

  PijGij \73:71 (P[73], \P72:71 , G[73], \G72:71 , \P73:71 , \G73:71 );

  wire \P73:63 , \G73:63 ;

  PijGij \73:63 (\P73:71 , \P70:63 , \G73:71 , \G70:63 , \P73:63 , \G73:63 );

  wire \G73:-1 ;

  Gij \73:-1 (\P73:63 , \G73:63 , \G62:-1 , \G73:-1 );

  Sum s74(\G73:-1 , A[74], B[74], S[74]);

  wire \P74:73 , \G74:73 ;

  PijGij \74:73 (P[74], P[73], G[74], G[73], \P74:73 , \G74:73 );

  wire \P74:71 , \G74:71 ;

  PijGij \74:71 (\P74:73 , \P72:71 , \G74:73 , \G72:71 , \P74:71 , \G74:71 );

  wire \P74:63 , \G74:63 ;

  PijGij \74:63 (\P74:71 , \P70:63 , \G74:71 , \G70:63 , \P74:63 , \G74:63 );

  wire \G74:-1 ;

  Gij \74:-1 (\P74:63 , \G74:63 , \G62:-1 , \G74:-1 );

  Sum s75(\G74:-1 , A[75], B[75], S[75]);

  wire \P75:71 , \G75:71 ;

  PijGij \75:71 (P[75], \P74:71 , G[75], \G74:71 , \P75:71 , \G75:71 );

  wire \P75:63 , \G75:63 ;

  PijGij \75:63 (\P75:71 , \P70:63 , \G75:71 , \G70:63 , \P75:63 , \G75:63 );

  wire \G75:-1 ;

  Gij \75:-1 (\P75:63 , \G75:63 , \G62:-1 , \G75:-1 );

  Sum s76(\G75:-1 , A[76], B[76], S[76]);

  wire \P76:75 , \G76:75 ;

  PijGij \76:75 (P[76], P[75], G[76], G[75], \P76:75 , \G76:75 );

  wire \P76:71 , \G76:71 ;

  PijGij \76:71 (\P76:75 , \P74:71 , \G76:75 , \G74:71 , \P76:71 , \G76:71 );

  wire \P76:63 , \G76:63 ;

  PijGij \76:63 (\P76:71 , \P70:63 , \G76:71 , \G70:63 , \P76:63 , \G76:63 );

  wire \G76:-1 ;

  Gij \76:-1 (\P76:63 , \G76:63 , \G62:-1 , \G76:-1 );

  Sum s77(\G76:-1 , A[77], B[77], S[77]);

  wire \P77:75 , \G77:75 ;

  PijGij \77:75 (P[77], \P76:75 , G[77], \G76:75 , \P77:75 , \G77:75 );

  wire \P77:71 , \G77:71 ;

  PijGij \77:71 (\P77:75 , \P74:71 , \G77:75 , \G74:71 , \P77:71 , \G77:71 );

  wire \P77:63 , \G77:63 ;

  PijGij \77:63 (\P77:71 , \P70:63 , \G77:71 , \G70:63 , \P77:63 , \G77:63 );

  wire \G77:-1 ;

  Gij \77:-1 (\P77:63 , \G77:63 , \G62:-1 , \G77:-1 );

  Sum s78(\G77:-1 , A[78], B[78], S[78]);

  wire \P78:77 , \G78:77 ;

  PijGij \78:77 (P[78], P[77], G[78], G[77], \P78:77 , \G78:77 );

  wire \P78:75 , \G78:75 ;

  PijGij \78:75 (\P78:77 , \P76:75 , \G78:77 , \G76:75 , \P78:75 , \G78:75 );

  wire \P78:71 , \G78:71 ;

  PijGij \78:71 (\P78:75 , \P74:71 , \G78:75 , \G74:71 , \P78:71 , \G78:71 );

  wire \P78:63 , \G78:63 ;

  PijGij \78:63 (\P78:71 , \P70:63 , \G78:71 , \G70:63 , \P78:63 , \G78:63 );

  wire \G78:-1 ;

  Gij \78:-1 (\P78:63 , \G78:63 , \G62:-1 , \G78:-1 );

  Sum s79(\G78:-1 , A[79], B[79], S[79]);

  wire \P79:63 , \G79:63 ;

  PijGij \79:63 (P[79], \P78:63 , G[79], \G78:63 , \P79:63 , \G79:63 );

  wire \G79:-1 ;

  Gij \79:-1 (\P79:63 , \G79:63 , \G62:-1 , \G79:-1 );

  Sum s80(\G79:-1 , A[80], B[80], S[80]);

  wire \P80:79 , \G80:79 ;

  PijGij \80:79 (P[80], P[79], G[80], G[79], \P80:79 , \G80:79 );

  wire \P80:63 , \G80:63 ;

  PijGij \80:63 (\P80:79 , \P78:63 , \G80:79 , \G78:63 , \P80:63 , \G80:63 );

  wire \G80:-1 ;

  Gij \80:-1 (\P80:63 , \G80:63 , \G62:-1 , \G80:-1 );

  Sum s81(\G80:-1 , A[81], B[81], S[81]);

  wire \P81:79 , \G81:79 ;

  PijGij \81:79 (P[81], \P80:79 , G[81], \G80:79 , \P81:79 , \G81:79 );

  wire \P81:63 , \G81:63 ;

  PijGij \81:63 (\P81:79 , \P78:63 , \G81:79 , \G78:63 , \P81:63 , \G81:63 );

  wire \G81:-1 ;

  Gij \81:-1 (\P81:63 , \G81:63 , \G62:-1 , \G81:-1 );

  Sum s82(\G81:-1 , A[82], B[82], S[82]);

  wire \P82:81 , \G82:81 ;

  PijGij \82:81 (P[82], P[81], G[82], G[81], \P82:81 , \G82:81 );

  wire \P82:79 , \G82:79 ;

  PijGij \82:79 (\P82:81 , \P80:79 , \G82:81 , \G80:79 , \P82:79 , \G82:79 );

  wire \P82:63 , \G82:63 ;

  PijGij \82:63 (\P82:79 , \P78:63 , \G82:79 , \G78:63 , \P82:63 , \G82:63 );

  wire \G82:-1 ;

  Gij \82:-1 (\P82:63 , \G82:63 , \G62:-1 , \G82:-1 );

  Sum s83(\G82:-1 , A[83], B[83], S[83]);

  wire \P83:79 , \G83:79 ;

  PijGij \83:79 (P[83], \P82:79 , G[83], \G82:79 , \P83:79 , \G83:79 );

  wire \P83:63 , \G83:63 ;

  PijGij \83:63 (\P83:79 , \P78:63 , \G83:79 , \G78:63 , \P83:63 , \G83:63 );

  wire \G83:-1 ;

  Gij \83:-1 (\P83:63 , \G83:63 , \G62:-1 , \G83:-1 );

  Sum s84(\G83:-1 , A[84], B[84], S[84]);

  wire \P84:83 , \G84:83 ;

  PijGij \84:83 (P[84], P[83], G[84], G[83], \P84:83 , \G84:83 );

  wire \P84:79 , \G84:79 ;

  PijGij \84:79 (\P84:83 , \P82:79 , \G84:83 , \G82:79 , \P84:79 , \G84:79 );

  wire \P84:63 , \G84:63 ;

  PijGij \84:63 (\P84:79 , \P78:63 , \G84:79 , \G78:63 , \P84:63 , \G84:63 );

  wire \G84:-1 ;

  Gij \84:-1 (\P84:63 , \G84:63 , \G62:-1 , \G84:-1 );

  Sum s85(\G84:-1 , A[85], B[85], S[85]);

  wire \P85:83 , \G85:83 ;

  PijGij \85:83 (P[85], \P84:83 , G[85], \G84:83 , \P85:83 , \G85:83 );

  wire \P85:79 , \G85:79 ;

  PijGij \85:79 (\P85:83 , \P82:79 , \G85:83 , \G82:79 , \P85:79 , \G85:79 );

  wire \P85:63 , \G85:63 ;

  PijGij \85:63 (\P85:79 , \P78:63 , \G85:79 , \G78:63 , \P85:63 , \G85:63 );

  wire \G85:-1 ;

  Gij \85:-1 (\P85:63 , \G85:63 , \G62:-1 , \G85:-1 );

  Sum s86(\G85:-1 , A[86], B[86], S[86]);

  wire \P86:85 , \G86:85 ;

  PijGij \86:85 (P[86], P[85], G[86], G[85], \P86:85 , \G86:85 );

  wire \P86:83 , \G86:83 ;

  PijGij \86:83 (\P86:85 , \P84:83 , \G86:85 , \G84:83 , \P86:83 , \G86:83 );

  wire \P86:79 , \G86:79 ;

  PijGij \86:79 (\P86:83 , \P82:79 , \G86:83 , \G82:79 , \P86:79 , \G86:79 );

  wire \P86:63 , \G86:63 ;

  PijGij \86:63 (\P86:79 , \P78:63 , \G86:79 , \G78:63 , \P86:63 , \G86:63 );

  wire \G86:-1 ;

  Gij \86:-1 (\P86:63 , \G86:63 , \G62:-1 , \G86:-1 );

  Sum s87(\G86:-1 , A[87], B[87], S[87]);

  wire \P87:79 , \G87:79 ;

  PijGij \87:79 (P[87], \P86:79 , G[87], \G86:79 , \P87:79 , \G87:79 );

  wire \P87:63 , \G87:63 ;

  PijGij \87:63 (\P87:79 , \P78:63 , \G87:79 , \G78:63 , \P87:63 , \G87:63 );

  wire \G87:-1 ;

  Gij \87:-1 (\P87:63 , \G87:63 , \G62:-1 , \G87:-1 );

  Sum s88(\G87:-1 , A[88], B[88], S[88]);

  wire \P88:87 , \G88:87 ;

  PijGij \88:87 (P[88], P[87], G[88], G[87], \P88:87 , \G88:87 );

  wire \P88:79 , \G88:79 ;

  PijGij \88:79 (\P88:87 , \P86:79 , \G88:87 , \G86:79 , \P88:79 , \G88:79 );

  wire \P88:63 , \G88:63 ;

  PijGij \88:63 (\P88:79 , \P78:63 , \G88:79 , \G78:63 , \P88:63 , \G88:63 );

  wire \G88:-1 ;

  Gij \88:-1 (\P88:63 , \G88:63 , \G62:-1 , \G88:-1 );

  Sum s89(\G88:-1 , A[89], B[89], S[89]);

  wire \P89:87 , \G89:87 ;

  PijGij \89:87 (P[89], \P88:87 , G[89], \G88:87 , \P89:87 , \G89:87 );

  wire \P89:79 , \G89:79 ;

  PijGij \89:79 (\P89:87 , \P86:79 , \G89:87 , \G86:79 , \P89:79 , \G89:79 );

  wire \P89:63 , \G89:63 ;

  PijGij \89:63 (\P89:79 , \P78:63 , \G89:79 , \G78:63 , \P89:63 , \G89:63 );

  wire \G89:-1 ;

  Gij \89:-1 (\P89:63 , \G89:63 , \G62:-1 , \G89:-1 );

  Sum s90(\G89:-1 , A[90], B[90], S[90]);

  wire \P90:89 , \G90:89 ;

  PijGij \90:89 (P[90], P[89], G[90], G[89], \P90:89 , \G90:89 );

  wire \P90:87 , \G90:87 ;

  PijGij \90:87 (\P90:89 , \P88:87 , \G90:89 , \G88:87 , \P90:87 , \G90:87 );

  wire \P90:79 , \G90:79 ;

  PijGij \90:79 (\P90:87 , \P86:79 , \G90:87 , \G86:79 , \P90:79 , \G90:79 );

  wire \P90:63 , \G90:63 ;

  PijGij \90:63 (\P90:79 , \P78:63 , \G90:79 , \G78:63 , \P90:63 , \G90:63 );

  wire \G90:-1 ;

  Gij \90:-1 (\P90:63 , \G90:63 , \G62:-1 , \G90:-1 );

  Sum s91(\G90:-1 , A[91], B[91], S[91]);

  wire \P91:87 , \G91:87 ;

  PijGij \91:87 (P[91], \P90:87 , G[91], \G90:87 , \P91:87 , \G91:87 );

  wire \P91:79 , \G91:79 ;

  PijGij \91:79 (\P91:87 , \P86:79 , \G91:87 , \G86:79 , \P91:79 , \G91:79 );

  wire \P91:63 , \G91:63 ;

  PijGij \91:63 (\P91:79 , \P78:63 , \G91:79 , \G78:63 , \P91:63 , \G91:63 );

  wire \G91:-1 ;

  Gij \91:-1 (\P91:63 , \G91:63 , \G62:-1 , \G91:-1 );

  Sum s92(\G91:-1 , A[92], B[92], S[92]);

  wire \P92:91 , \G92:91 ;

  PijGij \92:91 (P[92], P[91], G[92], G[91], \P92:91 , \G92:91 );

  wire \P92:87 , \G92:87 ;

  PijGij \92:87 (\P92:91 , \P90:87 , \G92:91 , \G90:87 , \P92:87 , \G92:87 );

  wire \P92:79 , \G92:79 ;

  PijGij \92:79 (\P92:87 , \P86:79 , \G92:87 , \G86:79 , \P92:79 , \G92:79 );

  wire \P92:63 , \G92:63 ;

  PijGij \92:63 (\P92:79 , \P78:63 , \G92:79 , \G78:63 , \P92:63 , \G92:63 );

  wire \G92:-1 ;

  Gij \92:-1 (\P92:63 , \G92:63 , \G62:-1 , \G92:-1 );

  Sum s93(\G92:-1 , A[93], B[93], S[93]);

  wire \P93:91 , \G93:91 ;

  PijGij \93:91 (P[93], \P92:91 , G[93], \G92:91 , \P93:91 , \G93:91 );

  wire \P93:87 , \G93:87 ;

  PijGij \93:87 (\P93:91 , \P90:87 , \G93:91 , \G90:87 , \P93:87 , \G93:87 );

  wire \P93:79 , \G93:79 ;

  PijGij \93:79 (\P93:87 , \P86:79 , \G93:87 , \G86:79 , \P93:79 , \G93:79 );

  wire \P93:63 , \G93:63 ;

  PijGij \93:63 (\P93:79 , \P78:63 , \G93:79 , \G78:63 , \P93:63 , \G93:63 );

  wire \G93:-1 ;

  Gij \93:-1 (\P93:63 , \G93:63 , \G62:-1 , \G93:-1 );

  Sum s94(\G93:-1 , A[94], B[94], S[94]);

  wire \P94:93 , \G94:93 ;

  PijGij \94:93 (P[94], P[93], G[94], G[93], \P94:93 , \G94:93 );

  wire \P94:91 , \G94:91 ;

  PijGij \94:91 (\P94:93 , \P92:91 , \G94:93 , \G92:91 , \P94:91 , \G94:91 );

  wire \P94:87 , \G94:87 ;

  PijGij \94:87 (\P94:91 , \P90:87 , \G94:91 , \G90:87 , \P94:87 , \G94:87 );

  wire \P94:79 , \G94:79 ;

  PijGij \94:79 (\P94:87 , \P86:79 , \G94:87 , \G86:79 , \P94:79 , \G94:79 );

  wire \P94:63 , \G94:63 ;

  PijGij \94:63 (\P94:79 , \P78:63 , \G94:79 , \G78:63 , \P94:63 , \G94:63 );

  wire \G94:-1 ;

  Gij \94:-1 (\P94:63 , \G94:63 , \G62:-1 , \G94:-1 );

  Sum s95(\G94:-1 , A[95], B[95], S[95]);

  wire \P95:63 , \G95:63 ;

  PijGij \95:63 (P[95], \P94:63 , G[95], \G94:63 , \P95:63 , \G95:63 );

  wire \G95:-1 ;

  Gij \95:-1 (\P95:63 , \G95:63 , \G62:-1 , \G95:-1 );

  Sum s96(\G95:-1 , A[96], B[96], S[96]);

  wire \P96:95 , \G96:95 ;

  PijGij \96:95 (P[96], P[95], G[96], G[95], \P96:95 , \G96:95 );

  wire \P96:63 , \G96:63 ;

  PijGij \96:63 (\P96:95 , \P94:63 , \G96:95 , \G94:63 , \P96:63 , \G96:63 );

  wire \G96:-1 ;

  Gij \96:-1 (\P96:63 , \G96:63 , \G62:-1 , \G96:-1 );

  Sum s97(\G96:-1 , A[97], B[97], S[97]);

  wire \P97:95 , \G97:95 ;

  PijGij \97:95 (P[97], \P96:95 , G[97], \G96:95 , \P97:95 , \G97:95 );

  wire \P97:63 , \G97:63 ;

  PijGij \97:63 (\P97:95 , \P94:63 , \G97:95 , \G94:63 , \P97:63 , \G97:63 );

  wire \G97:-1 ;

  Gij \97:-1 (\P97:63 , \G97:63 , \G62:-1 , \G97:-1 );

  Sum s98(\G97:-1 , A[98], B[98], S[98]);

  wire \P98:97 , \G98:97 ;

  PijGij \98:97 (P[98], P[97], G[98], G[97], \P98:97 , \G98:97 );

  wire \P98:95 , \G98:95 ;

  PijGij \98:95 (\P98:97 , \P96:95 , \G98:97 , \G96:95 , \P98:95 , \G98:95 );

  wire \P98:63 , \G98:63 ;

  PijGij \98:63 (\P98:95 , \P94:63 , \G98:95 , \G94:63 , \P98:63 , \G98:63 );

  wire \G98:-1 ;

  Gij \98:-1 (\P98:63 , \G98:63 , \G62:-1 , \G98:-1 );

  Sum s99(\G98:-1 , A[99], B[99], S[99]);

  wire \P99:95 , \G99:95 ;

  PijGij \99:95 (P[99], \P98:95 , G[99], \G98:95 , \P99:95 , \G99:95 );

  wire \P99:63 , \G99:63 ;

  PijGij \99:63 (\P99:95 , \P94:63 , \G99:95 , \G94:63 , \P99:63 , \G99:63 );

  wire \G99:-1 ;

  Gij \99:-1 (\P99:63 , \G99:63 , \G62:-1 , \G99:-1 );

  Sum s100(\G99:-1 , A[100], B[100], S[100]);

  wire \P100:99 , \G100:99 ;

  PijGij \100:99 (P[100], P[99], G[100], G[99], \P100:99 , \G100:99 );

  wire \P100:95 , \G100:95 ;

  PijGij \100:95 (\P100:99 , \P98:95 , \G100:99 , \G98:95 , \P100:95 , \G100:95 );

  wire \P100:63 , \G100:63 ;

  PijGij \100:63 (\P100:95 , \P94:63 , \G100:95 , \G94:63 , \P100:63 , \G100:63 );

  wire \G100:-1 ;

  Gij \100:-1 (\P100:63 , \G100:63 , \G62:-1 , \G100:-1 );

  Sum s101(\G100:-1 , A[101], B[101], S[101]);

  wire \P101:99 , \G101:99 ;

  PijGij \101:99 (P[101], \P100:99 , G[101], \G100:99 , \P101:99 , \G101:99 );

  wire \P101:95 , \G101:95 ;

  PijGij \101:95 (\P101:99 , \P98:95 , \G101:99 , \G98:95 , \P101:95 , \G101:95 );

  wire \P101:63 , \G101:63 ;

  PijGij \101:63 (\P101:95 , \P94:63 , \G101:95 , \G94:63 , \P101:63 , \G101:63 );

  wire \G101:-1 ;

  Gij \101:-1 (\P101:63 , \G101:63 , \G62:-1 , \G101:-1 );

  Sum s102(\G101:-1 , A[102], B[102], S[102]);

  wire \P102:101 , \G102:101 ;

  PijGij \102:101 (P[102], P[101], G[102], G[101], \P102:101 , \G102:101 );

  wire \P102:99 , \G102:99 ;

  PijGij \102:99 (\P102:101 , \P100:99 , \G102:101 , \G100:99 , \P102:99 , \G102:99 );

  wire \P102:95 , \G102:95 ;

  PijGij \102:95 (\P102:99 , \P98:95 , \G102:99 , \G98:95 , \P102:95 , \G102:95 );

  wire \P102:63 , \G102:63 ;

  PijGij \102:63 (\P102:95 , \P94:63 , \G102:95 , \G94:63 , \P102:63 , \G102:63 );

  wire \G102:-1 ;

  Gij \102:-1 (\P102:63 , \G102:63 , \G62:-1 , \G102:-1 );

  Sum s103(\G102:-1 , A[103], B[103], S[103]);

  wire \P103:95 , \G103:95 ;

  PijGij \103:95 (P[103], \P102:95 , G[103], \G102:95 , \P103:95 , \G103:95 );

  wire \P103:63 , \G103:63 ;

  PijGij \103:63 (\P103:95 , \P94:63 , \G103:95 , \G94:63 , \P103:63 , \G103:63 );

  wire \G103:-1 ;

  Gij \103:-1 (\P103:63 , \G103:63 , \G62:-1 , \G103:-1 );

  Sum s104(\G103:-1 , A[104], B[104], S[104]);

  wire \P104:103 , \G104:103 ;

  PijGij \104:103 (P[104], P[103], G[104], G[103], \P104:103 , \G104:103 );

  wire \P104:95 , \G104:95 ;

  PijGij \104:95 (\P104:103 , \P102:95 , \G104:103 , \G102:95 , \P104:95 , \G104:95 );

  wire \P104:63 , \G104:63 ;

  PijGij \104:63 (\P104:95 , \P94:63 , \G104:95 , \G94:63 , \P104:63 , \G104:63 );

  wire \G104:-1 ;

  Gij \104:-1 (\P104:63 , \G104:63 , \G62:-1 , \G104:-1 );

  Sum s105(\G104:-1 , A[105], B[105], S[105]);

  wire \P105:103 , \G105:103 ;

  PijGij \105:103 (P[105], \P104:103 , G[105], \G104:103 , \P105:103 , \G105:103 );

  wire \P105:95 , \G105:95 ;

  PijGij \105:95 (\P105:103 , \P102:95 , \G105:103 , \G102:95 , \P105:95 , \G105:95 );

  wire \P105:63 , \G105:63 ;

  PijGij \105:63 (\P105:95 , \P94:63 , \G105:95 , \G94:63 , \P105:63 , \G105:63 );

  wire \G105:-1 ;

  Gij \105:-1 (\P105:63 , \G105:63 , \G62:-1 , \G105:-1 );

  Sum s106(\G105:-1 , A[106], B[106], S[106]);

  wire \P106:105 , \G106:105 ;

  PijGij \106:105 (P[106], P[105], G[106], G[105], \P106:105 , \G106:105 );

  wire \P106:103 , \G106:103 ;

  PijGij \106:103 (\P106:105 , \P104:103 , \G106:105 , \G104:103 , \P106:103 , \G106:103 );

  wire \P106:95 , \G106:95 ;

  PijGij \106:95 (\P106:103 , \P102:95 , \G106:103 , \G102:95 , \P106:95 , \G106:95 );

  wire \P106:63 , \G106:63 ;

  PijGij \106:63 (\P106:95 , \P94:63 , \G106:95 , \G94:63 , \P106:63 , \G106:63 );

  wire \G106:-1 ;

  Gij \106:-1 (\P106:63 , \G106:63 , \G62:-1 , \G106:-1 );

  Sum s107(\G106:-1 , A[107], B[107], S[107]);

  wire \P107:103 , \G107:103 ;

  PijGij \107:103 (P[107], \P106:103 , G[107], \G106:103 , \P107:103 , \G107:103 );

  wire \P107:95 , \G107:95 ;

  PijGij \107:95 (\P107:103 , \P102:95 , \G107:103 , \G102:95 , \P107:95 , \G107:95 );

  wire \P107:63 , \G107:63 ;

  PijGij \107:63 (\P107:95 , \P94:63 , \G107:95 , \G94:63 , \P107:63 , \G107:63 );

  wire \G107:-1 ;

  Gij \107:-1 (\P107:63 , \G107:63 , \G62:-1 , \G107:-1 );

  Sum s108(\G107:-1 , A[108], B[108], S[108]);

  wire \P108:107 , \G108:107 ;

  PijGij \108:107 (P[108], P[107], G[108], G[107], \P108:107 , \G108:107 );

  wire \P108:103 , \G108:103 ;

  PijGij \108:103 (\P108:107 , \P106:103 , \G108:107 , \G106:103 , \P108:103 , \G108:103 );

  wire \P108:95 , \G108:95 ;

  PijGij \108:95 (\P108:103 , \P102:95 , \G108:103 , \G102:95 , \P108:95 , \G108:95 );

  wire \P108:63 , \G108:63 ;

  PijGij \108:63 (\P108:95 , \P94:63 , \G108:95 , \G94:63 , \P108:63 , \G108:63 );

  wire \G108:-1 ;

  Gij \108:-1 (\P108:63 , \G108:63 , \G62:-1 , \G108:-1 );

  Sum s109(\G108:-1 , A[109], B[109], S[109]);

  wire \P109:107 , \G109:107 ;

  PijGij \109:107 (P[109], \P108:107 , G[109], \G108:107 , \P109:107 , \G109:107 );

  wire \P109:103 , \G109:103 ;

  PijGij \109:103 (\P109:107 , \P106:103 , \G109:107 , \G106:103 , \P109:103 , \G109:103 );

  wire \P109:95 , \G109:95 ;

  PijGij \109:95 (\P109:103 , \P102:95 , \G109:103 , \G102:95 , \P109:95 , \G109:95 );

  wire \P109:63 , \G109:63 ;

  PijGij \109:63 (\P109:95 , \P94:63 , \G109:95 , \G94:63 , \P109:63 , \G109:63 );

  wire \G109:-1 ;

  Gij \109:-1 (\P109:63 , \G109:63 , \G62:-1 , \G109:-1 );

  Sum s110(\G109:-1 , A[110], B[110], S[110]);

  wire \P110:109 , \G110:109 ;

  PijGij \110:109 (P[110], P[109], G[110], G[109], \P110:109 , \G110:109 );

  wire \P110:107 , \G110:107 ;

  PijGij \110:107 (\P110:109 , \P108:107 , \G110:109 , \G108:107 , \P110:107 , \G110:107 );

  wire \P110:103 , \G110:103 ;

  PijGij \110:103 (\P110:107 , \P106:103 , \G110:107 , \G106:103 , \P110:103 , \G110:103 );

  wire \P110:95 , \G110:95 ;

  PijGij \110:95 (\P110:103 , \P102:95 , \G110:103 , \G102:95 , \P110:95 , \G110:95 );

  wire \P110:63 , \G110:63 ;

  PijGij \110:63 (\P110:95 , \P94:63 , \G110:95 , \G94:63 , \P110:63 , \G110:63 );

  wire \G110:-1 ;

  Gij \110:-1 (\P110:63 , \G110:63 , \G62:-1 , \G110:-1 );

  Sum s111(\G110:-1 , A[111], B[111], S[111]);

  wire \P111:95 , \G111:95 ;

  PijGij \111:95 (P[111], \P110:95 , G[111], \G110:95 , \P111:95 , \G111:95 );

  wire \P111:63 , \G111:63 ;

  PijGij \111:63 (\P111:95 , \P94:63 , \G111:95 , \G94:63 , \P111:63 , \G111:63 );

  wire \G111:-1 ;

  Gij \111:-1 (\P111:63 , \G111:63 , \G62:-1 , \G111:-1 );

  Sum s112(\G111:-1 , A[112], B[112], S[112]);

  assign Cout = (\G111:-1 & A[112]) | (\G111:-1 & B[112]) | (A[112] & B[112]);

endmodule
